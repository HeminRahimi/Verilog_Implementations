module Cross_mult (clk, r_cross, P0_prime, P1_prime, Q0_prime, Q1_prime, F0, F1);

        input clk;
        input [7 : 0] r_cross;
        input [14 : 0] P0_prime, P1_prime, Q0_prime, Q1_prime;
        output [7 : 0] F0, F1;

        assign  {a_0, b_0, c_0, d_0, ab_0, ac_0, ad_0, bc_0, bd_0, cd_0, abc_0, abd_0, acd_0, bcd_0, abcd_0} = P0_prime;
        assign  {a_1, b_1, c_1, d_1, ab_1, ac_1, ad_1, bc_1, bd_1, cd_1, abc_1, abd_1, acd_1, bcd_1, abcd_1} = P1_prime;
        
        assign {e_0, f_0, g_0, h_0, ef_0, eg_0, eh_0, fg_0, fh_0, gh_0, efg_0, efh_0, egh_0, fgh_0, efgh_0} = Q0_prime;
        assign {e_1, f_1, g_1, h_1, ef_1, eg_1, eh_1, fg_1, fh_1, gh_1, efg_1, efh_1, egh_1, fgh_1, efgh_1} = Q1_prime;

        assign f0_00 = h_0 ^ gh_0 ^ f_0 ^ fg_0 ^ e_0 ^ eg_0 ^ ef_0 ^ efg_0 ^ efgh_0 ^ d_0 ^ d_0 & h_0 ^ d_0 & g_0 ^ d_0 & gh_0 ^ d_0 & f_0 ^ d_0 & fh_0 ^ d_0 & fg_0 ^ d_0 & eh_0 ^ d_0 & eg_0 ^ d_0 & efgh_0 ^ c_0 & h_0 ^ c_0 & fh_0 ^ c_0 & fgh_0 ^ c_0 & eh_0 ^ c_0 & ef_0 ^ c_0 & efh_0 ^ c_0 & efg_0 ^ cd_0 & gh_0 ^ cd_0 & fh_0 ^ cd_0 & fgh_0 ^ cd_0 & efh_0 ^ b_0 & h_0 ^ b_0 & g_0 ^ b_0 & gh_0 ^ b_0 & f_0 ^ b_0 & fh_0 ^ b_0 & fg_0 ^ b_0 & fgh_0 ^ b_0 & eh_0 ^ b_0 & efg_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & h_0 ^ bd_0 & g_0 ^ bd_0 & fg_0 ^ bd_0 & eh_0 ^ bd_0 & eg_0 ^ bd_0 & egh_0 ^ bd_0 & efh_0 ^ bd_0 & efgh_0 ^ bc_0 ^ bc_0 & g_0 ^ bc_0 & f_0 ^ bc_0 & fh_0 ^ bc_0 & eh_0 ^ bc_0 & egh_0 ^ bc_0 & efg_0 ^ bcd_0 ^ bcd_0 & h_0 ^ bcd_0 & g_0 ^ bcd_0 & gh_0 ^ bcd_0 & f_0 ^ bcd_0 & fg_0 ^ bcd_0 & eh_0 ^ bcd_0 & ef_0 ^ bcd_0 & efh_0 ^ a_0 & gh_0 ^ a_0 & f_0 ^ a_0 & fh_0 ^ a_0 & fgh_0 ^ a_0 & eg_0 ^ a_0 & ef_0 ^ a_0 & efh_0 ^ a_0 & efg_0 ^ a_0 & efgh_0 ^ ad_0 & h_0 ^ ad_0 & gh_0 ^ ad_0 & f_0 ^ ad_0 & fh_0 ^ ad_0 & fg_0 ^ ad_0 & fgh_0 ^ ad_0 & e_0 ^ ad_0 & efgh_0 ^ ac_0 ^ ac_0 & f_0 ^ ac_0 & fh_0 ^ ac_0 & fgh_0 ^ ac_0 & e_0 ^ ac_0 & egh_0 ^ ac_0 & ef_0 ^ ac_0 & efg_0 ^ ac_0 & efgh_0 ^ acd_0 & h_0 ^ acd_0 & g_0 ^ acd_0 & f_0 ^ acd_0 & fh_0 ^ acd_0 & fgh_0 ^ acd_0 & eh_0 ^ acd_0 & eg_0 ^ acd_0 & ef_0 ^ acd_0 & efh_0 ^ ab_0 ^ ab_0 & f_0 ^ ab_0 & fg_0 ^ ab_0 & fgh_0 ^ ab_0 & e_0 ^ ab_0 & eg_0 ^ ab_0 & egh_0 ^ ab_0 & ef_0 ^ ab_0 & efgh_0 ^ abd_0 & h_0 ^ abd_0 & fh_0 ^ abd_0 & fg_0 ^ abd_0 & eh_0 ^ abd_0 & egh_0 ^ abd_0 & efg_0 ^ abd_0 & efgh_0 ^ abc_0 ^ abc_0 & g_0 ^ abc_0 & gh_0 ^ abc_0 & fg_0 ^ abc_0 & fgh_0 ^ abc_0 & e_0 ^ abc_0 & eh_0 ^ abc_0 & efh_0 ^ abcd_0 & gh_0 ^ abcd_0 & f_0 ^ abcd_0 & fg_0 ^ abcd_0 & fgh_0 ^ abcd_0 & eg_0 ^ abcd_0 & ef_0 ^ abcd_0 & efh_0 ;
        assign f0_01 = d_0 & h_1 ^ d_0 & g_1 ^ d_0 & gh_1 ^ d_0 & f_1 ^ d_0 & fh_1 ^ d_0 & fg_1 ^ d_0 & eh_1 ^ d_0 & eg_1 ^ d_0 & efgh_1 ^ c_0 & h_1 ^ c_0 & fh_1 ^ c_0 & fgh_1 ^ c_0 & eh_1 ^ c_0 & ef_1 ^ c_0 & efh_1 ^ c_0 & efg_1 ^ cd_0 & gh_1 ^ cd_0 & fh_1 ^ cd_0 & fgh_1 ^ cd_0 & efh_1 ^ b_0 & h_1 ^ b_0 & g_1 ^ b_0 & gh_1 ^ b_0 & f_1 ^ b_0 & fh_1 ^ b_0 & fg_1 ^ b_0 & fgh_1 ^ b_0 & eh_1 ^ b_0 & efg_1 ^ b_0 & efgh_1 ^ bd_0 & h_1 ^ bd_0 & g_1 ^ bd_0 & fg_1 ^ bd_0 & eh_1 ^ bd_0 & eg_1 ^ bd_0 & egh_1 ^ bd_0 & efh_1 ^ bd_0 & efgh_1 ^ bc_0 & g_1 ^ bc_0 & f_1 ^ bc_0 & fh_1 ^ bc_0 & eh_1 ^ bc_0 & egh_1 ^ bc_0 & efg_1 ^ bcd_0 & h_1 ^ bcd_0 & g_1 ^ bcd_0 & gh_1 ^ bcd_0 & f_1 ^ bcd_0 & fg_1 ^ bcd_0 & eh_1 ^ bcd_0 & ef_1 ^ bcd_0 & efh_1 ^ a_0 & gh_1 ^ a_0 & f_1 ^ a_0 & fh_1 ^ a_0 & fgh_1 ^ a_0 & eg_1 ^ a_0 & ef_1 ^ a_0 & efh_1 ^ a_0 & efg_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & gh_1 ^ ad_0 & f_1 ^ ad_0 & fh_1 ^ ad_0 & fg_1 ^ ad_0 & fgh_1 ^ ad_0 & e_1 ^ ad_0 & efgh_1 ^ ac_0 & f_1 ^ ac_0 & fh_1 ^ ac_0 & fgh_1 ^ ac_0 & e_1 ^ ac_0 & egh_1 ^ ac_0 & ef_1 ^ ac_0 & efg_1 ^ ac_0 & efgh_1 ^ acd_0 & h_1 ^ acd_0 & g_1 ^ acd_0 & f_1 ^ acd_0 & fh_1 ^ acd_0 & fgh_1 ^ acd_0 & eh_1 ^ acd_0 & eg_1 ^ acd_0 & ef_1 ^ acd_0 & efh_1 ^ ab_0 & f_1 ^ ab_0 & fg_1 ^ ab_0 & fgh_1 ^ ab_0 & e_1 ^ ab_0 & eg_1 ^ ab_0 & egh_1 ^ ab_0 & ef_1 ^ ab_0 & efgh_1 ^ abd_0 & h_1 ^ abd_0 & fh_1 ^ abd_0 & fg_1 ^ abd_0 & eh_1 ^ abd_0 & egh_1 ^ abd_0 & efg_1 ^ abd_0 & efgh_1 ^ abc_0 & g_1 ^ abc_0 & gh_1 ^ abc_0 & fg_1 ^ abc_0 & fgh_1 ^ abc_0 & e_1 ^ abc_0 & eh_1 ^ abc_0 & efh_1 ^ abcd_0 & gh_1 ^ abcd_0 & f_1 ^ abcd_0 & fg_1 ^ abcd_0 & fgh_1 ^ abcd_0 & eg_1 ^ abcd_0 & ef_1 ^ abcd_0 & efh_1 ;
        assign f0_10 = d_1 & h_0 ^ d_1 & g_0 ^ d_1 & gh_0 ^ d_1 & f_0 ^ d_1 & fh_0 ^ d_1 & fg_0 ^ d_1 & eh_0 ^ d_1 & eg_0 ^ d_1 & efgh_0 ^ c_1 & h_0 ^ c_1 & fh_0 ^ c_1 & fgh_0 ^ c_1 & eh_0 ^ c_1 & ef_0 ^ c_1 & efh_0 ^ c_1 & efg_0 ^ cd_1 & gh_0 ^ cd_1 & fh_0 ^ cd_1 & fgh_0 ^ cd_1 & efh_0 ^ b_1 & h_0 ^ b_1 & g_0 ^ b_1 & gh_0 ^ b_1 & f_0 ^ b_1 & fh_0 ^ b_1 & fg_0 ^ b_1 & fgh_0 ^ b_1 & eh_0 ^ b_1 & efg_0 ^ b_1 & efgh_0 ^ bd_1 & h_0 ^ bd_1 & g_0 ^ bd_1 & fg_0 ^ bd_1 & eh_0 ^ bd_1 & eg_0 ^ bd_1 & egh_0 ^ bd_1 & efh_0 ^ bd_1 & efgh_0 ^ bc_1 & g_0 ^ bc_1 & f_0 ^ bc_1 & fh_0 ^ bc_1 & eh_0 ^ bc_1 & egh_0 ^ bc_1 & efg_0 ^ bcd_1 & h_0 ^ bcd_1 & g_0 ^ bcd_1 & gh_0 ^ bcd_1 & f_0 ^ bcd_1 & fg_0 ^ bcd_1 & eh_0 ^ bcd_1 & ef_0 ^ bcd_1 & efh_0 ^ a_1 & gh_0 ^ a_1 & f_0 ^ a_1 & fh_0 ^ a_1 & fgh_0 ^ a_1 & eg_0 ^ a_1 & ef_0 ^ a_1 & efh_0 ^ a_1 & efg_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & gh_0 ^ ad_1 & f_0 ^ ad_1 & fh_0 ^ ad_1 & fg_0 ^ ad_1 & fgh_0 ^ ad_1 & e_0 ^ ad_1 & efgh_0 ^ ac_1 & f_0 ^ ac_1 & fh_0 ^ ac_1 & fgh_0 ^ ac_1 & e_0 ^ ac_1 & egh_0 ^ ac_1 & ef_0 ^ ac_1 & efg_0 ^ ac_1 & efgh_0 ^ acd_1 & h_0 ^ acd_1 & g_0 ^ acd_1 & f_0 ^ acd_1 & fh_0 ^ acd_1 & fgh_0 ^ acd_1 & eh_0 ^ acd_1 & eg_0 ^ acd_1 & ef_0 ^ acd_1 & efh_0 ^ ab_1 & f_0 ^ ab_1 & fg_0 ^ ab_1 & fgh_0 ^ ab_1 & e_0 ^ ab_1 & eg_0 ^ ab_1 & egh_0 ^ ab_1 & ef_0 ^ ab_1 & efgh_0 ^ abd_1 & h_0 ^ abd_1 & fh_0 ^ abd_1 & fg_0 ^ abd_1 & eh_0 ^ abd_1 & egh_0 ^ abd_1 & efg_0 ^ abd_1 & efgh_0 ^ abc_1 & g_0 ^ abc_1 & gh_0 ^ abc_1 & fg_0 ^ abc_1 & fgh_0 ^ abc_1 & e_0 ^ abc_1 & eh_0 ^ abc_1 & efh_0 ^ abcd_1 & gh_0 ^ abcd_1 & f_0 ^ abcd_1 & fg_0 ^ abcd_1 & fgh_0 ^ abcd_1 & eg_0 ^ abcd_1 & ef_0 ^ abcd_1 & efh_0 ;
        assign f0_11 = h_1 ^ gh_1 ^ f_1 ^ fg_1 ^ e_1 ^ eg_1 ^ ef_1 ^ efg_1 ^ efgh_1 ^ d_1 ^ d_1 & h_1 ^ d_1 & g_1 ^ d_1 & gh_1 ^ d_1 & f_1 ^ d_1 & fh_1 ^ d_1 & fg_1 ^ d_1 & eh_1 ^ d_1 & eg_1 ^ d_1 & efgh_1 ^ c_1 & h_1 ^ c_1 & fh_1 ^ c_1 & fgh_1 ^ c_1 & eh_1 ^ c_1 & ef_1 ^ c_1 & efh_1 ^ c_1 & efg_1 ^ cd_1 & gh_1 ^ cd_1 & fh_1 ^ cd_1 & fgh_1 ^ cd_1 & efh_1 ^ b_1 & h_1 ^ b_1 & g_1 ^ b_1 & gh_1 ^ b_1 & f_1 ^ b_1 & fh_1 ^ b_1 & fg_1 ^ b_1 & fgh_1 ^ b_1 & eh_1 ^ b_1 & efg_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & h_1 ^ bd_1 & g_1 ^ bd_1 & fg_1 ^ bd_1 & eh_1 ^ bd_1 & eg_1 ^ bd_1 & egh_1 ^ bd_1 & efh_1 ^ bd_1 & efgh_1 ^ bc_1 ^ bc_1 & g_1 ^ bc_1 & f_1 ^ bc_1 & fh_1 ^ bc_1 & eh_1 ^ bc_1 & egh_1 ^ bc_1 & efg_1 ^ bcd_1 ^ bcd_1 & h_1 ^ bcd_1 & g_1 ^ bcd_1 & gh_1 ^ bcd_1 & f_1 ^ bcd_1 & fg_1 ^ bcd_1 & eh_1 ^ bcd_1 & ef_1 ^ bcd_1 & efh_1 ^ a_1 & gh_1 ^ a_1 & f_1 ^ a_1 & fh_1 ^ a_1 & fgh_1 ^ a_1 & eg_1 ^ a_1 & ef_1 ^ a_1 & efh_1 ^ a_1 & efg_1 ^ a_1 & efgh_1 ^ ad_1 & h_1 ^ ad_1 & gh_1 ^ ad_1 & f_1 ^ ad_1 & fh_1 ^ ad_1 & fg_1 ^ ad_1 & fgh_1 ^ ad_1 & e_1 ^ ad_1 & efgh_1 ^ ac_1 ^ ac_1 & f_1 ^ ac_1 & fh_1 ^ ac_1 & fgh_1 ^ ac_1 & e_1 ^ ac_1 & egh_1 ^ ac_1 & ef_1 ^ ac_1 & efg_1 ^ ac_1 & efgh_1 ^ acd_1 & h_1 ^ acd_1 & g_1 ^ acd_1 & f_1 ^ acd_1 & fh_1 ^ acd_1 & fgh_1 ^ acd_1 & eh_1 ^ acd_1 & eg_1 ^ acd_1 & ef_1 ^ acd_1 & efh_1 ^ ab_1 ^ ab_1 & f_1 ^ ab_1 & fg_1 ^ ab_1 & fgh_1 ^ ab_1 & e_1 ^ ab_1 & eg_1 ^ ab_1 & egh_1 ^ ab_1 & ef_1 ^ ab_1 & efgh_1 ^ abd_1 & h_1 ^ abd_1 & fh_1 ^ abd_1 & fg_1 ^ abd_1 & eh_1 ^ abd_1 & egh_1 ^ abd_1 & efg_1 ^ abd_1 & efgh_1 ^ abc_1 ^ abc_1 & g_1 ^ abc_1 & gh_1 ^ abc_1 & fg_1 ^ abc_1 & fgh_1 ^ abc_1 & e_1 ^ abc_1 & eh_1 ^ abc_1 & efh_1 ^ abcd_1 & gh_1 ^ abcd_1 & f_1 ^ abcd_1 & fg_1 ^ abcd_1 & fgh_1 ^ abcd_1 & eg_1 ^ abcd_1 & ef_1 ^ abcd_1 & efh_1 ;
        wire f0_00_reg;
        Register # (1) inst_inner_f0_00 (f0_00, clk, f0_00_reg);
        wire f0_01_reg;
        Register # (1) inst_cross_f0_01 (f0_01 ^ r_cross[0], clk, f0_01_reg);
        wire f0_10_reg;
        Register # (1) inst_cross_f0_10 (f0_10 ^ r_cross[0], clk, f0_10_reg);
        wire f0_11_reg;
        Register # (1) inst_inner_f0_11 (f0_11, clk, f0_11_reg);
        
        assign f1_00 = h_0 ^ gh_0 ^ fh_0 ^ e_0 ^ eh_0 ^ eg_0 ^ egh_0 ^ ef_0 ^ efh_0 ^ efg_0 ^ d_0 & h_0 ^ d_0 & g_0 ^ d_0 & gh_0 ^ d_0 & fg_0 ^ d_0 & eh_0 ^ d_0 & eg_0 ^ d_0 & egh_0 ^ d_0 & ef_0 ^ d_0 & efgh_0 ^ c_0 & eg_0 ^ c_0 & ef_0 ^ c_0 & efg_0 ^ cd_0 ^ cd_0 & h_0 ^ cd_0 & gh_0 ^ cd_0 & fh_0 ^ cd_0 & fgh_0 ^ cd_0 & eh_0 ^ cd_0 & eg_0 ^ cd_0 & ef_0 ^ cd_0 & efh_0 ^ b_0 ^ b_0 & gh_0 ^ b_0 & f_0 ^ b_0 & fgh_0 ^ b_0 & eg_0 ^ b_0 & egh_0 ^ b_0 & ef_0 ^ b_0 & efh_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & h_0 ^ bd_0 & fgh_0 ^ bd_0 & e_0 ^ bd_0 & eh_0 ^ bd_0 & egh_0 ^ bd_0 & efg_0 ^ bd_0 & efgh_0 ^ bc_0 & g_0 ^ bc_0 & gh_0 ^ bc_0 & fh_0 ^ bc_0 & fg_0 ^ bc_0 & e_0 ^ bc_0 & eg_0 ^ bc_0 & egh_0 ^ bc_0 & efg_0 ^ bc_0 & efgh_0 ^ bcd_0 & h_0 ^ bcd_0 & gh_0 ^ bcd_0 & fh_0 ^ bcd_0 & fg_0 ^ bcd_0 & e_0 ^ bcd_0 & eg_0 ^ bcd_0 & egh_0 ^ bcd_0 & efh_0 ^ bcd_0 & efg_0 ^ a_0 ^ a_0 & h_0 ^ a_0 & g_0 ^ a_0 & f_0 ^ a_0 & fh_0 ^ a_0 & e_0 ^ a_0 & eg_0 ^ a_0 & efgh_0 ^ ad_0 & h_0 ^ ad_0 & g_0 ^ ad_0 & gh_0 ^ ad_0 & fg_0 ^ ad_0 & fgh_0 ^ ad_0 & e_0 ^ ad_0 & eg_0 ^ ad_0 & egh_0 ^ ad_0 & ef_0 ^ ad_0 & efh_0 ^ ad_0 & efgh_0 ^ ac_0 & h_0 ^ ac_0 & f_0 ^ ac_0 & fg_0 ^ ac_0 & e_0 ^ ac_0 & eg_0 ^ ac_0 & egh_0 ^ ac_0 & ef_0 ^ ac_0 & efh_0 ^ acd_0 & h_0 ^ acd_0 & g_0 ^ acd_0 & f_0 ^ acd_0 & fgh_0 ^ acd_0 & e_0 ^ acd_0 & eh_0 ^ acd_0 & eg_0 ^ acd_0 & ef_0 ^ acd_0 & efh_0 ^ ab_0 & h_0 ^ ab_0 & f_0 ^ ab_0 & fg_0 ^ ab_0 & fgh_0 ^ ab_0 & e_0 ^ ab_0 & egh_0 ^ ab_0 & efh_0 ^ abd_0 & h_0 ^ abd_0 & g_0 ^ abd_0 & f_0 ^ abd_0 & fgh_0 ^ abd_0 & e_0 ^ abd_0 & egh_0 ^ abd_0 & ef_0 ^ abd_0 & efh_0 ^ abd_0 & efg_0 ^ abd_0 & efgh_0 ^ abc_0 ^ abc_0 & gh_0 ^ abc_0 & fh_0 ^ abc_0 & fgh_0 ^ abc_0 & eh_0 ^ abc_0 & efh_0 ^ abc_0 & efg_0 ^ abc_0 & efgh_0 ^ abcd_0 & h_0 ^ abcd_0 & f_0 ^ abcd_0 & fgh_0 ^ abcd_0 & eg_0 ^ abcd_0 & egh_0 ;
        assign f1_01 = d_0 & h_1 ^ d_0 & g_1 ^ d_0 & gh_1 ^ d_0 & fg_1 ^ d_0 & eh_1 ^ d_0 & eg_1 ^ d_0 & egh_1 ^ d_0 & ef_1 ^ d_0 & efgh_1 ^ c_0 & eg_1 ^ c_0 & ef_1 ^ c_0 & efg_1 ^ cd_0 & h_1 ^ cd_0 & gh_1 ^ cd_0 & fh_1 ^ cd_0 & fgh_1 ^ cd_0 & eh_1 ^ cd_0 & eg_1 ^ cd_0 & ef_1 ^ cd_0 & efh_1 ^ b_0 & gh_1 ^ b_0 & f_1 ^ b_0 & fgh_1 ^ b_0 & eg_1 ^ b_0 & egh_1 ^ b_0 & ef_1 ^ b_0 & efh_1 ^ b_0 & efgh_1 ^ bd_0 & h_1 ^ bd_0 & fgh_1 ^ bd_0 & e_1 ^ bd_0 & eh_1 ^ bd_0 & egh_1 ^ bd_0 & efg_1 ^ bd_0 & efgh_1 ^ bc_0 & g_1 ^ bc_0 & gh_1 ^ bc_0 & fh_1 ^ bc_0 & fg_1 ^ bc_0 & e_1 ^ bc_0 & eg_1 ^ bc_0 & egh_1 ^ bc_0 & efg_1 ^ bc_0 & efgh_1 ^ bcd_0 & h_1 ^ bcd_0 & gh_1 ^ bcd_0 & fh_1 ^ bcd_0 & fg_1 ^ bcd_0 & e_1 ^ bcd_0 & eg_1 ^ bcd_0 & egh_1 ^ bcd_0 & efh_1 ^ bcd_0 & efg_1 ^ a_0 & h_1 ^ a_0 & g_1 ^ a_0 & f_1 ^ a_0 & fh_1 ^ a_0 & e_1 ^ a_0 & eg_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & g_1 ^ ad_0 & gh_1 ^ ad_0 & fg_1 ^ ad_0 & fgh_1 ^ ad_0 & e_1 ^ ad_0 & eg_1 ^ ad_0 & egh_1 ^ ad_0 & ef_1 ^ ad_0 & efh_1 ^ ad_0 & efgh_1 ^ ac_0 & h_1 ^ ac_0 & f_1 ^ ac_0 & fg_1 ^ ac_0 & e_1 ^ ac_0 & eg_1 ^ ac_0 & egh_1 ^ ac_0 & ef_1 ^ ac_0 & efh_1 ^ acd_0 & h_1 ^ acd_0 & g_1 ^ acd_0 & f_1 ^ acd_0 & fgh_1 ^ acd_0 & e_1 ^ acd_0 & eh_1 ^ acd_0 & eg_1 ^ acd_0 & ef_1 ^ acd_0 & efh_1 ^ ab_0 & h_1 ^ ab_0 & f_1 ^ ab_0 & fg_1 ^ ab_0 & fgh_1 ^ ab_0 & e_1 ^ ab_0 & egh_1 ^ ab_0 & efh_1 ^ abd_0 & h_1 ^ abd_0 & g_1 ^ abd_0 & f_1 ^ abd_0 & fgh_1 ^ abd_0 & e_1 ^ abd_0 & egh_1 ^ abd_0 & ef_1 ^ abd_0 & efh_1 ^ abd_0 & efg_1 ^ abd_0 & efgh_1 ^ abc_0 & gh_1 ^ abc_0 & fh_1 ^ abc_0 & fgh_1 ^ abc_0 & eh_1 ^ abc_0 & efh_1 ^ abc_0 & efg_1 ^ abc_0 & efgh_1 ^ abcd_0 & h_1 ^ abcd_0 & f_1 ^ abcd_0 & fgh_1 ^ abcd_0 & eg_1 ^ abcd_0 & egh_1 ;
        assign f1_10 = d_1 & h_0 ^ d_1 & g_0 ^ d_1 & gh_0 ^ d_1 & fg_0 ^ d_1 & eh_0 ^ d_1 & eg_0 ^ d_1 & egh_0 ^ d_1 & ef_0 ^ d_1 & efgh_0 ^ c_1 & eg_0 ^ c_1 & ef_0 ^ c_1 & efg_0 ^ cd_1 & h_0 ^ cd_1 & gh_0 ^ cd_1 & fh_0 ^ cd_1 & fgh_0 ^ cd_1 & eh_0 ^ cd_1 & eg_0 ^ cd_1 & ef_0 ^ cd_1 & efh_0 ^ b_1 & gh_0 ^ b_1 & f_0 ^ b_1 & fgh_0 ^ b_1 & eg_0 ^ b_1 & egh_0 ^ b_1 & ef_0 ^ b_1 & efh_0 ^ b_1 & efgh_0 ^ bd_1 & h_0 ^ bd_1 & fgh_0 ^ bd_1 & e_0 ^ bd_1 & eh_0 ^ bd_1 & egh_0 ^ bd_1 & efg_0 ^ bd_1 & efgh_0 ^ bc_1 & g_0 ^ bc_1 & gh_0 ^ bc_1 & fh_0 ^ bc_1 & fg_0 ^ bc_1 & e_0 ^ bc_1 & eg_0 ^ bc_1 & egh_0 ^ bc_1 & efg_0 ^ bc_1 & efgh_0 ^ bcd_1 & h_0 ^ bcd_1 & gh_0 ^ bcd_1 & fh_0 ^ bcd_1 & fg_0 ^ bcd_1 & e_0 ^ bcd_1 & eg_0 ^ bcd_1 & egh_0 ^ bcd_1 & efh_0 ^ bcd_1 & efg_0 ^ a_1 & h_0 ^ a_1 & g_0 ^ a_1 & f_0 ^ a_1 & fh_0 ^ a_1 & e_0 ^ a_1 & eg_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & g_0 ^ ad_1 & gh_0 ^ ad_1 & fg_0 ^ ad_1 & fgh_0 ^ ad_1 & e_0 ^ ad_1 & eg_0 ^ ad_1 & egh_0 ^ ad_1 & ef_0 ^ ad_1 & efh_0 ^ ad_1 & efgh_0 ^ ac_1 & h_0 ^ ac_1 & f_0 ^ ac_1 & fg_0 ^ ac_1 & e_0 ^ ac_1 & eg_0 ^ ac_1 & egh_0 ^ ac_1 & ef_0 ^ ac_1 & efh_0 ^ acd_1 & h_0 ^ acd_1 & g_0 ^ acd_1 & f_0 ^ acd_1 & fgh_0 ^ acd_1 & e_0 ^ acd_1 & eh_0 ^ acd_1 & eg_0 ^ acd_1 & ef_0 ^ acd_1 & efh_0 ^ ab_1 & h_0 ^ ab_1 & f_0 ^ ab_1 & fg_0 ^ ab_1 & fgh_0 ^ ab_1 & e_0 ^ ab_1 & egh_0 ^ ab_1 & efh_0 ^ abd_1 & h_0 ^ abd_1 & g_0 ^ abd_1 & f_0 ^ abd_1 & fgh_0 ^ abd_1 & e_0 ^ abd_1 & egh_0 ^ abd_1 & ef_0 ^ abd_1 & efh_0 ^ abd_1 & efg_0 ^ abd_1 & efgh_0 ^ abc_1 & gh_0 ^ abc_1 & fh_0 ^ abc_1 & fgh_0 ^ abc_1 & eh_0 ^ abc_1 & efh_0 ^ abc_1 & efg_0 ^ abc_1 & efgh_0 ^ abcd_1 & h_0 ^ abcd_1 & f_0 ^ abcd_1 & fgh_0 ^ abcd_1 & eg_0 ^ abcd_1 & egh_0 ;
        assign f1_11 = h_1 ^ gh_1 ^ fh_1 ^ e_1 ^ eh_1 ^ eg_1 ^ egh_1 ^ ef_1 ^ efh_1 ^ efg_1 ^ d_1 & h_1 ^ d_1 & g_1 ^ d_1 & gh_1 ^ d_1 & fg_1 ^ d_1 & eh_1 ^ d_1 & eg_1 ^ d_1 & egh_1 ^ d_1 & ef_1 ^ d_1 & efgh_1 ^ c_1 & eg_1 ^ c_1 & ef_1 ^ c_1 & efg_1 ^ cd_1 ^ cd_1 & h_1 ^ cd_1 & gh_1 ^ cd_1 & fh_1 ^ cd_1 & fgh_1 ^ cd_1 & eh_1 ^ cd_1 & eg_1 ^ cd_1 & ef_1 ^ cd_1 & efh_1 ^ b_1 ^ b_1 & gh_1 ^ b_1 & f_1 ^ b_1 & fgh_1 ^ b_1 & eg_1 ^ b_1 & egh_1 ^ b_1 & ef_1 ^ b_1 & efh_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & h_1 ^ bd_1 & fgh_1 ^ bd_1 & e_1 ^ bd_1 & eh_1 ^ bd_1 & egh_1 ^ bd_1 & efg_1 ^ bd_1 & efgh_1 ^ bc_1 & g_1 ^ bc_1 & gh_1 ^ bc_1 & fh_1 ^ bc_1 & fg_1 ^ bc_1 & e_1 ^ bc_1 & eg_1 ^ bc_1 & egh_1 ^ bc_1 & efg_1 ^ bc_1 & efgh_1 ^ bcd_1 & h_1 ^ bcd_1 & gh_1 ^ bcd_1 & fh_1 ^ bcd_1 & fg_1 ^ bcd_1 & e_1 ^ bcd_1 & eg_1 ^ bcd_1 & egh_1 ^ bcd_1 & efh_1 ^ bcd_1 & efg_1 ^ a_1 ^ a_1 & h_1 ^ a_1 & g_1 ^ a_1 & f_1 ^ a_1 & fh_1 ^ a_1 & e_1 ^ a_1 & eg_1 ^ a_1 & efgh_1 ^ ad_1 & h_1 ^ ad_1 & g_1 ^ ad_1 & gh_1 ^ ad_1 & fg_1 ^ ad_1 & fgh_1 ^ ad_1 & e_1 ^ ad_1 & eg_1 ^ ad_1 & egh_1 ^ ad_1 & ef_1 ^ ad_1 & efh_1 ^ ad_1 & efgh_1 ^ ac_1 & h_1 ^ ac_1 & f_1 ^ ac_1 & fg_1 ^ ac_1 & e_1 ^ ac_1 & eg_1 ^ ac_1 & egh_1 ^ ac_1 & ef_1 ^ ac_1 & efh_1 ^ acd_1 & h_1 ^ acd_1 & g_1 ^ acd_1 & f_1 ^ acd_1 & fgh_1 ^ acd_1 & e_1 ^ acd_1 & eh_1 ^ acd_1 & eg_1 ^ acd_1 & ef_1 ^ acd_1 & efh_1 ^ ab_1 & h_1 ^ ab_1 & f_1 ^ ab_1 & fg_1 ^ ab_1 & fgh_1 ^ ab_1 & e_1 ^ ab_1 & egh_1 ^ ab_1 & efh_1 ^ abd_1 & h_1 ^ abd_1 & g_1 ^ abd_1 & f_1 ^ abd_1 & fgh_1 ^ abd_1 & e_1 ^ abd_1 & egh_1 ^ abd_1 & ef_1 ^ abd_1 & efh_1 ^ abd_1 & efg_1 ^ abd_1 & efgh_1 ^ abc_1 ^ abc_1 & gh_1 ^ abc_1 & fh_1 ^ abc_1 & fgh_1 ^ abc_1 & eh_1 ^ abc_1 & efh_1 ^ abc_1 & efg_1 ^ abc_1 & efgh_1 ^ abcd_1 & h_1 ^ abcd_1 & f_1 ^ abcd_1 & fgh_1 ^ abcd_1 & eg_1 ^ abcd_1 & egh_1 ;
        wire f1_00_reg;
        Register # (1) inst_inner_f1_00 (f1_00, clk, f1_00_reg);
        wire f1_01_reg;
        Register # (1) inst_cross_f1_01 (f1_01 ^ r_cross[1], clk, f1_01_reg);
        wire f1_10_reg;
        Register # (1) inst_cross_f1_10 (f1_10 ^ r_cross[1], clk, f1_10_reg);
        wire f1_11_reg;
        Register # (1) inst_inner_f1_11 (f1_11, clk, f1_11_reg);
        ///////////////
        
        assign f2_00 = h_0 ^ g_0 ^ fh_0 ^ eh_0 ^ egh_0 ^ ef_0 ^ efh_0 ^ d_0 & h_0 ^ d_0 & g_0 ^ d_0 & gh_0 ^ d_0 & fh_0 ^ d_0 & fg_0 ^ d_0 & e_0 ^ d_0 & eh_0 ^ d_0 & eg_0 ^ d_0 & egh_0 ^ d_0 & ef_0 ^ d_0 & efh_0 ^ d_0 & efg_0 ^ d_0 & efgh_0 ^ c_0 ^ c_0 & h_0 ^ c_0 & gh_0 ^ c_0 & fh_0 ^ c_0 & fg_0 ^ c_0 & fgh_0 ^ c_0 & eh_0 ^ c_0 & eg_0 ^ c_0 & egh_0 ^ c_0 & efh_0 ^ c_0 & efg_0 ^ c_0 & efgh_0 ^ cd_0 & h_0 ^ cd_0 & g_0 ^ cd_0 & f_0 ^ cd_0 & fgh_0 ^ cd_0 & e_0 ^ cd_0 & efg_0 ^ cd_0 & efgh_0 ^ b_0 & h_0 ^ b_0 & gh_0 ^ b_0 & fg_0 ^ b_0 & eh_0 ^ b_0 & egh_0 ^ b_0 & ef_0 ^ b_0 & efg_0 ^ b_0 & efgh_0 ^ bd_0 & h_0 ^ bd_0 & gh_0 ^ bd_0 & fh_0 ^ bd_0 & e_0 ^ bd_0 & eh_0 ^ bd_0 & egh_0 ^ bd_0 & ef_0 ^ bd_0 & efg_0 ^ bd_0 & efgh_0 ^ bc_0 ^ bc_0 & g_0 ^ bc_0 & gh_0 ^ bc_0 & e_0 ^ bc_0 & eh_0 ^ bc_0 & ef_0 ^ bc_0 & efgh_0 ^ bcd_0 & f_0 ^ bcd_0 & fh_0 ^ bcd_0 & fg_0 ^ bcd_0 & fgh_0 ^ bcd_0 & e_0 ^ bcd_0 & eg_0 ^ bcd_0 & efh_0 ^ a_0 ^ a_0 & h_0 ^ a_0 & gh_0 ^ a_0 & fh_0 ^ a_0 & fg_0 ^ a_0 & fgh_0 ^ a_0 & eh_0 ^ a_0 & eg_0 ^ a_0 & ef_0 ^ a_0 & efh_0 ^ a_0 & efgh_0 ^ ad_0 ^ ad_0 & h_0 ^ ad_0 & g_0 ^ ad_0 & fh_0 ^ ad_0 & fg_0 ^ ad_0 & fgh_0 ^ ad_0 & eh_0 ^ ad_0 & egh_0 ^ ad_0 & ef_0 ^ ad_0 & efh_0 ^ ad_0 & efgh_0 ^ ac_0 & h_0 ^ ac_0 & g_0 ^ ac_0 & fg_0 ^ ac_0 & fgh_0 ^ ac_0 & eh_0 ^ ac_0 & eg_0 ^ ac_0 & egh_0 ^ ac_0 & efh_0 ^ acd_0 & g_0 ^ acd_0 & f_0 ^ acd_0 & fg_0 ^ acd_0 & fgh_0 ^ acd_0 & eh_0 ^ acd_0 & egh_0 ^ acd_0 & efg_0 ^ ab_0 ^ ab_0 & h_0 ^ ab_0 & f_0 ^ ab_0 & fg_0 ^ ab_0 & fgh_0 ^ ab_0 & eg_0 ^ ab_0 & egh_0 ^ ab_0 & efg_0 ^ abd_0 ^ abd_0 & gh_0 ^ abd_0 & f_0 ^ abd_0 & fg_0 ^ abd_0 & eg_0 ^ abd_0 & egh_0 ^ abd_0 & ef_0 ^ abd_0 & efh_0 ^ abd_0 & efg_0 ^ abd_0 & efgh_0 ^ abc_0 & g_0 ^ abc_0 & f_0 ^ abc_0 & fh_0 ^ abc_0 & e_0 ^ abc_0 & eh_0 ^ abc_0 & eg_0 ^ abc_0 & egh_0 ^ abc_0 & ef_0 ^ abc_0 & efh_0 ^ abc_0 & efgh_0 ^ abcd_0 ^ abcd_0 & h_0 ^ abcd_0 & g_0 ^ abcd_0 & gh_0 ^ abcd_0 & fh_0 ^ abcd_0 & e_0 ^ abcd_0 & egh_0 ^ abcd_0 & ef_0 ^ abcd_0 & efh_0 ^ abcd_0 & efg_0 ;
        assign f2_01 = d_0 & h_1 ^ d_0 & g_1 ^ d_0 & gh_1 ^ d_0 & fh_1 ^ d_0 & fg_1 ^ d_0 & e_1 ^ d_0 & eh_1 ^ d_0 & eg_1 ^ d_0 & egh_1 ^ d_0 & ef_1 ^ d_0 & efh_1 ^ d_0 & efg_1 ^ d_0 & efgh_1 ^ c_0 & h_1 ^ c_0 & gh_1 ^ c_0 & fh_1 ^ c_0 & fg_1 ^ c_0 & fgh_1 ^ c_0 & eh_1 ^ c_0 & eg_1 ^ c_0 & egh_1 ^ c_0 & efh_1 ^ c_0 & efg_1 ^ c_0 & efgh_1 ^ cd_0 & h_1 ^ cd_0 & g_1 ^ cd_0 & f_1 ^ cd_0 & fgh_1 ^ cd_0 & e_1 ^ cd_0 & efg_1 ^ cd_0 & efgh_1 ^ b_0 & h_1 ^ b_0 & gh_1 ^ b_0 & fg_1 ^ b_0 & eh_1 ^ b_0 & egh_1 ^ b_0 & ef_1 ^ b_0 & efg_1 ^ b_0 & efgh_1 ^ bd_0 & h_1 ^ bd_0 & gh_1 ^ bd_0 & fh_1 ^ bd_0 & e_1 ^ bd_0 & eh_1 ^ bd_0 & egh_1 ^ bd_0 & ef_1 ^ bd_0 & efg_1 ^ bd_0 & efgh_1 ^ bc_0 & g_1 ^ bc_0 & gh_1 ^ bc_0 & e_1 ^ bc_0 & eh_1 ^ bc_0 & ef_1 ^ bc_0 & efgh_1 ^ bcd_0 & f_1 ^ bcd_0 & fh_1 ^ bcd_0 & fg_1 ^ bcd_0 & fgh_1 ^ bcd_0 & e_1 ^ bcd_0 & eg_1 ^ bcd_0 & efh_1 ^ a_0 & h_1 ^ a_0 & gh_1 ^ a_0 & fh_1 ^ a_0 & fg_1 ^ a_0 & fgh_1 ^ a_0 & eh_1 ^ a_0 & eg_1 ^ a_0 & ef_1 ^ a_0 & efh_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & g_1 ^ ad_0 & fh_1 ^ ad_0 & fg_1 ^ ad_0 & fgh_1 ^ ad_0 & eh_1 ^ ad_0 & egh_1 ^ ad_0 & ef_1 ^ ad_0 & efh_1 ^ ad_0 & efgh_1 ^ ac_0 & h_1 ^ ac_0 & g_1 ^ ac_0 & fg_1 ^ ac_0 & fgh_1 ^ ac_0 & eh_1 ^ ac_0 & eg_1 ^ ac_0 & egh_1 ^ ac_0 & efh_1 ^ acd_0 & g_1 ^ acd_0 & f_1 ^ acd_0 & fg_1 ^ acd_0 & fgh_1 ^ acd_0 & eh_1 ^ acd_0 & egh_1 ^ acd_0 & efg_1 ^ ab_0 & h_1 ^ ab_0 & f_1 ^ ab_0 & fg_1 ^ ab_0 & fgh_1 ^ ab_0 & eg_1 ^ ab_0 & egh_1 ^ ab_0 & efg_1 ^ abd_0 & gh_1 ^ abd_0 & f_1 ^ abd_0 & fg_1 ^ abd_0 & eg_1 ^ abd_0 & egh_1 ^ abd_0 & ef_1 ^ abd_0 & efh_1 ^ abd_0 & efg_1 ^ abd_0 & efgh_1 ^ abc_0 & g_1 ^ abc_0 & f_1 ^ abc_0 & fh_1 ^ abc_0 & e_1 ^ abc_0 & eh_1 ^ abc_0 & eg_1 ^ abc_0 & egh_1 ^ abc_0 & ef_1 ^ abc_0 & efh_1 ^ abc_0 & efgh_1 ^ abcd_0 & h_1 ^ abcd_0 & g_1 ^ abcd_0 & gh_1 ^ abcd_0 & fh_1 ^ abcd_0 & e_1 ^ abcd_0 & egh_1 ^ abcd_0 & ef_1 ^ abcd_0 & efh_1 ^ abcd_0 & efg_1 ;
        assign f2_10 = d_1 & h_0 ^ d_1 & g_0 ^ d_1 & gh_0 ^ d_1 & fh_0 ^ d_1 & fg_0 ^ d_1 & e_0 ^ d_1 & eh_0 ^ d_1 & eg_0 ^ d_1 & egh_0 ^ d_1 & ef_0 ^ d_1 & efh_0 ^ d_1 & efg_0 ^ d_1 & efgh_0 ^ c_1 & h_0 ^ c_1 & gh_0 ^ c_1 & fh_0 ^ c_1 & fg_0 ^ c_1 & fgh_0 ^ c_1 & eh_0 ^ c_1 & eg_0 ^ c_1 & egh_0 ^ c_1 & efh_0 ^ c_1 & efg_0 ^ c_1 & efgh_0 ^ cd_1 & h_0 ^ cd_1 & g_0 ^ cd_1 & f_0 ^ cd_1 & fgh_0 ^ cd_1 & e_0 ^ cd_1 & efg_0 ^ cd_1 & efgh_0 ^ b_1 & h_0 ^ b_1 & gh_0 ^ b_1 & fg_0 ^ b_1 & eh_0 ^ b_1 & egh_0 ^ b_1 & ef_0 ^ b_1 & efg_0 ^ b_1 & efgh_0 ^ bd_1 & h_0 ^ bd_1 & gh_0 ^ bd_1 & fh_0 ^ bd_1 & e_0 ^ bd_1 & eh_0 ^ bd_1 & egh_0 ^ bd_1 & ef_0 ^ bd_1 & efg_0 ^ bd_1 & efgh_0 ^ bc_1 & g_0 ^ bc_1 & gh_0 ^ bc_1 & e_0 ^ bc_1 & eh_0 ^ bc_1 & ef_0 ^ bc_1 & efgh_0 ^ bcd_1 & f_0 ^ bcd_1 & fh_0 ^ bcd_1 & fg_0 ^ bcd_1 & fgh_0 ^ bcd_1 & e_0 ^ bcd_1 & eg_0 ^ bcd_1 & efh_0 ^ a_1 & h_0 ^ a_1 & gh_0 ^ a_1 & fh_0 ^ a_1 & fg_0 ^ a_1 & fgh_0 ^ a_1 & eh_0 ^ a_1 & eg_0 ^ a_1 & ef_0 ^ a_1 & efh_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & g_0 ^ ad_1 & fh_0 ^ ad_1 & fg_0 ^ ad_1 & fgh_0 ^ ad_1 & eh_0 ^ ad_1 & egh_0 ^ ad_1 & ef_0 ^ ad_1 & efh_0 ^ ad_1 & efgh_0 ^ ac_1 & h_0 ^ ac_1 & g_0 ^ ac_1 & fg_0 ^ ac_1 & fgh_0 ^ ac_1 & eh_0 ^ ac_1 & eg_0 ^ ac_1 & egh_0 ^ ac_1 & efh_0 ^ acd_1 & g_0 ^ acd_1 & f_0 ^ acd_1 & fg_0 ^ acd_1 & fgh_0 ^ acd_1 & eh_0 ^ acd_1 & egh_0 ^ acd_1 & efg_0 ^ ab_1 & h_0 ^ ab_1 & f_0 ^ ab_1 & fg_0 ^ ab_1 & fgh_0 ^ ab_1 & eg_0 ^ ab_1 & egh_0 ^ ab_1 & efg_0 ^ abd_1 & gh_0 ^ abd_1 & f_0 ^ abd_1 & fg_0 ^ abd_1 & eg_0 ^ abd_1 & egh_0 ^ abd_1 & ef_0 ^ abd_1 & efh_0 ^ abd_1 & efg_0 ^ abd_1 & efgh_0 ^ abc_1 & g_0 ^ abc_1 & f_0 ^ abc_1 & fh_0 ^ abc_1 & e_0 ^ abc_1 & eh_0 ^ abc_1 & eg_0 ^ abc_1 & egh_0 ^ abc_1 & ef_0 ^ abc_1 & efh_0 ^ abc_1 & efgh_0 ^ abcd_1 & h_0 ^ abcd_1 & g_0 ^ abcd_1 & gh_0 ^ abcd_1 & fh_0 ^ abcd_1 & e_0 ^ abcd_1 & egh_0 ^ abcd_1 & ef_0 ^ abcd_1 & efh_0 ^ abcd_1 & efg_0 ;
        assign f2_11 = h_1 ^ g_1 ^ fh_1 ^ eh_1 ^ egh_1 ^ ef_1 ^ efh_1 ^ d_1 & h_1 ^ d_1 & g_1 ^ d_1 & gh_1 ^ d_1 & fh_1 ^ d_1 & fg_1 ^ d_1 & e_1 ^ d_1 & eh_1 ^ d_1 & eg_1 ^ d_1 & egh_1 ^ d_1 & ef_1 ^ d_1 & efh_1 ^ d_1 & efg_1 ^ d_1 & efgh_1 ^ c_1 ^ c_1 & h_1 ^ c_1 & gh_1 ^ c_1 & fh_1 ^ c_1 & fg_1 ^ c_1 & fgh_1 ^ c_1 & eh_1 ^ c_1 & eg_1 ^ c_1 & egh_1 ^ c_1 & efh_1 ^ c_1 & efg_1 ^ c_1 & efgh_1 ^ cd_1 & h_1 ^ cd_1 & g_1 ^ cd_1 & f_1 ^ cd_1 & fgh_1 ^ cd_1 & e_1 ^ cd_1 & efg_1 ^ cd_1 & efgh_1 ^ b_1 & h_1 ^ b_1 & gh_1 ^ b_1 & fg_1 ^ b_1 & eh_1 ^ b_1 & egh_1 ^ b_1 & ef_1 ^ b_1 & efg_1 ^ b_1 & efgh_1 ^ bd_1 & h_1 ^ bd_1 & gh_1 ^ bd_1 & fh_1 ^ bd_1 & e_1 ^ bd_1 & eh_1 ^ bd_1 & egh_1 ^ bd_1 & ef_1 ^ bd_1 & efg_1 ^ bd_1 & efgh_1 ^ bc_1 ^ bc_1 & g_1 ^ bc_1 & gh_1 ^ bc_1 & e_1 ^ bc_1 & eh_1 ^ bc_1 & ef_1 ^ bc_1 & efgh_1 ^ bcd_1 & f_1 ^ bcd_1 & fh_1 ^ bcd_1 & fg_1 ^ bcd_1 & fgh_1 ^ bcd_1 & e_1 ^ bcd_1 & eg_1 ^ bcd_1 & efh_1 ^ a_1 ^ a_1 & h_1 ^ a_1 & gh_1 ^ a_1 & fh_1 ^ a_1 & fg_1 ^ a_1 & fgh_1 ^ a_1 & eh_1 ^ a_1 & eg_1 ^ a_1 & ef_1 ^ a_1 & efh_1 ^ a_1 & efgh_1 ^ ad_1 ^ ad_1 & h_1 ^ ad_1 & g_1 ^ ad_1 & fh_1 ^ ad_1 & fg_1 ^ ad_1 & fgh_1 ^ ad_1 & eh_1 ^ ad_1 & egh_1 ^ ad_1 & ef_1 ^ ad_1 & efh_1 ^ ad_1 & efgh_1 ^ ac_1 & h_1 ^ ac_1 & g_1 ^ ac_1 & fg_1 ^ ac_1 & fgh_1 ^ ac_1 & eh_1 ^ ac_1 & eg_1 ^ ac_1 & egh_1 ^ ac_1 & efh_1 ^ acd_1 & g_1 ^ acd_1 & f_1 ^ acd_1 & fg_1 ^ acd_1 & fgh_1 ^ acd_1 & eh_1 ^ acd_1 & egh_1 ^ acd_1 & efg_1 ^ ab_1 ^ ab_1 & h_1 ^ ab_1 & f_1 ^ ab_1 & fg_1 ^ ab_1 & fgh_1 ^ ab_1 & eg_1 ^ ab_1 & egh_1 ^ ab_1 & efg_1 ^ abd_1 ^ abd_1 & gh_1 ^ abd_1 & f_1 ^ abd_1 & fg_1 ^ abd_1 & eg_1 ^ abd_1 & egh_1 ^ abd_1 & ef_1 ^ abd_1 & efh_1 ^ abd_1 & efg_1 ^ abd_1 & efgh_1 ^ abc_1 & g_1 ^ abc_1 & f_1 ^ abc_1 & fh_1 ^ abc_1 & e_1 ^ abc_1 & eh_1 ^ abc_1 & eg_1 ^ abc_1 & egh_1 ^ abc_1 & ef_1 ^ abc_1 & efh_1 ^ abc_1 & efgh_1 ^ abcd_1 ^ abcd_1 & h_1 ^ abcd_1 & g_1 ^ abcd_1 & gh_1 ^ abcd_1 & fh_1 ^ abcd_1 & e_1 ^ abcd_1 & egh_1 ^ abcd_1 & ef_1 ^ abcd_1 & efh_1 ^ abcd_1 & efg_1 ;
        wire f2_00_reg;
        Register # (1) inst_inner_f2_00 (f2_00, clk, f2_00_reg);
        wire f2_01_reg;
        Register # (1) inst_cross_f2_01 (f2_01 ^ r_cross[2], clk, f2_01_reg);
        wire f2_10_reg;
        Register # (1) inst_cross_f2_10 (f2_10 ^ r_cross[2], clk, f2_10_reg);
        wire f2_11_reg;
        Register # (1) inst_inner_f2_11 (f2_11, clk, f2_11_reg);
        ///////////////
        
        assign f3_00 = h_0 ^ fg_0 ^ eh_0 ^ egh_0 ^ ef_0 ^ efh_0 ^ efg_0 ^ efgh_0 ^ d_0 ^ d_0 & gh_0 ^ d_0 & fh_0 ^ d_0 & fgh_0 ^ d_0 & eh_0 ^ d_0 & eg_0 ^ d_0 & ef_0 ^ d_0 & efgh_0 ^ c_0 & gh_0 ^ c_0 & fg_0 ^ c_0 & fgh_0 ^ c_0 & ef_0 ^ c_0 & efg_0 ^ c_0 & efgh_0 ^ cd_0 ^ cd_0 & h_0 ^ cd_0 & f_0 ^ cd_0 & fg_0 ^ cd_0 & eg_0 ^ cd_0 & egh_0 ^ cd_0 & ef_0 ^ cd_0 & efh_0 ^ b_0 ^ b_0 & gh_0 ^ b_0 & fh_0 ^ b_0 & fg_0 ^ b_0 & e_0 ^ b_0 & eh_0 ^ b_0 & egh_0 ^ b_0 & efg_0 ^ bd_0 & h_0 ^ bd_0 & gh_0 ^ bd_0 & fh_0 ^ bd_0 & eh_0 ^ bd_0 & eg_0 ^ bd_0 & egh_0 ^ bd_0 & efgh_0 ^ bc_0 ^ bc_0 & g_0 ^ bc_0 & gh_0 ^ bc_0 & fh_0 ^ bc_0 & fgh_0 ^ bc_0 & e_0 ^ bc_0 & eg_0 ^ bc_0 & egh_0 ^ bc_0 & efh_0 ^ bc_0 & efg_0 ^ bc_0 & efgh_0 ^ bcd_0 & h_0 ^ bcd_0 & g_0 ^ bcd_0 & f_0 ^ bcd_0 & fh_0 ^ bcd_0 & fg_0 ^ bcd_0 & e_0 ^ bcd_0 & eh_0 ^ bcd_0 & ef_0 ^ bcd_0 & efg_0 ^ bcd_0 & efgh_0 ^ a_0 ^ a_0 & h_0 ^ a_0 & g_0 ^ a_0 & gh_0 ^ a_0 & fh_0 ^ a_0 & fg_0 ^ a_0 & e_0 ^ a_0 & eh_0 ^ a_0 & ef_0 ^ a_0 & efh_0 ^ a_0 & efg_0 ^ a_0 & efgh_0 ^ ad_0 & fh_0 ^ ad_0 & fg_0 ^ ad_0 & fgh_0 ^ ad_0 & e_0 ^ ad_0 & eg_0 ^ ad_0 & egh_0 ^ ad_0 & efgh_0 ^ ac_0 ^ ac_0 & f_0 ^ ac_0 & fg_0 ^ ac_0 & fgh_0 ^ ac_0 & e_0 ^ ac_0 & efh_0 ^ ac_0 & efgh_0 ^ acd_0 & g_0 ^ acd_0 & gh_0 ^ acd_0 & f_0 ^ acd_0 & fh_0 ^ acd_0 & fgh_0 ^ acd_0 & eh_0 ^ acd_0 & egh_0 ^ acd_0 & ef_0 ^ acd_0 & efg_0 ^ ab_0 ^ ab_0 & gh_0 ^ ab_0 & fh_0 ^ ab_0 & fg_0 ^ ab_0 & eh_0 ^ ab_0 & efh_0 ^ ab_0 & efgh_0 ^ abd_0 & g_0 ^ abd_0 & f_0 ^ abd_0 & fgh_0 ^ abd_0 & e_0 ^ abd_0 & eh_0 ^ abd_0 & eg_0 ^ abd_0 & efh_0 ^ abd_0 & efg_0 ^ abc_0 ^ abc_0 & h_0 ^ abc_0 & g_0 ^ abc_0 & gh_0 ^ abc_0 & fh_0 ^ abc_0 & fg_0 ^ abc_0 & e_0 ^ abc_0 & eh_0 ^ abc_0 & eg_0 ^ abc_0 & efh_0 ^ abc_0 & efg_0 ^ abc_0 & efgh_0 ^ abcd_0 ^ abcd_0 & h_0 ^ abcd_0 & f_0 ^ abcd_0 & fg_0 ^ abcd_0 & e_0 ^ abcd_0 & egh_0 ^ abcd_0 & ef_0 ^ abcd_0 & efh_0 ;
        assign f3_01 = d_0 & gh_1 ^ d_0 & fh_1 ^ d_0 & fgh_1 ^ d_0 & eh_1 ^ d_0 & eg_1 ^ d_0 & ef_1 ^ d_0 & efgh_1 ^ c_0 & gh_1 ^ c_0 & fg_1 ^ c_0 & fgh_1 ^ c_0 & ef_1 ^ c_0 & efg_1 ^ c_0 & efgh_1 ^ cd_0 & h_1 ^ cd_0 & f_1 ^ cd_0 & fg_1 ^ cd_0 & eg_1 ^ cd_0 & egh_1 ^ cd_0 & ef_1 ^ cd_0 & efh_1 ^ b_0 & gh_1 ^ b_0 & fh_1 ^ b_0 & fg_1 ^ b_0 & e_1 ^ b_0 & eh_1 ^ b_0 & egh_1 ^ b_0 & efg_1 ^ bd_0 & h_1 ^ bd_0 & gh_1 ^ bd_0 & fh_1 ^ bd_0 & eh_1 ^ bd_0 & eg_1 ^ bd_0 & egh_1 ^ bd_0 & efgh_1 ^ bc_0 & g_1 ^ bc_0 & gh_1 ^ bc_0 & fh_1 ^ bc_0 & fgh_1 ^ bc_0 & e_1 ^ bc_0 & eg_1 ^ bc_0 & egh_1 ^ bc_0 & efh_1 ^ bc_0 & efg_1 ^ bc_0 & efgh_1 ^ bcd_0 & h_1 ^ bcd_0 & g_1 ^ bcd_0 & f_1 ^ bcd_0 & fh_1 ^ bcd_0 & fg_1 ^ bcd_0 & e_1 ^ bcd_0 & eh_1 ^ bcd_0 & ef_1 ^ bcd_0 & efg_1 ^ bcd_0 & efgh_1 ^ a_0 & h_1 ^ a_0 & g_1 ^ a_0 & gh_1 ^ a_0 & fh_1 ^ a_0 & fg_1 ^ a_0 & e_1 ^ a_0 & eh_1 ^ a_0 & ef_1 ^ a_0 & efh_1 ^ a_0 & efg_1 ^ a_0 & efgh_1 ^ ad_0 & fh_1 ^ ad_0 & fg_1 ^ ad_0 & fgh_1 ^ ad_0 & e_1 ^ ad_0 & eg_1 ^ ad_0 & egh_1 ^ ad_0 & efgh_1 ^ ac_0 & f_1 ^ ac_0 & fg_1 ^ ac_0 & fgh_1 ^ ac_0 & e_1 ^ ac_0 & efh_1 ^ ac_0 & efgh_1 ^ acd_0 & g_1 ^ acd_0 & gh_1 ^ acd_0 & f_1 ^ acd_0 & fh_1 ^ acd_0 & fgh_1 ^ acd_0 & eh_1 ^ acd_0 & egh_1 ^ acd_0 & ef_1 ^ acd_0 & efg_1 ^ ab_0 & gh_1 ^ ab_0 & fh_1 ^ ab_0 & fg_1 ^ ab_0 & eh_1 ^ ab_0 & efh_1 ^ ab_0 & efgh_1 ^ abd_0 & g_1 ^ abd_0 & f_1 ^ abd_0 & fgh_1 ^ abd_0 & e_1 ^ abd_0 & eh_1 ^ abd_0 & eg_1 ^ abd_0 & efh_1 ^ abd_0 & efg_1 ^ abc_0 & h_1 ^ abc_0 & g_1 ^ abc_0 & gh_1 ^ abc_0 & fh_1 ^ abc_0 & fg_1 ^ abc_0 & e_1 ^ abc_0 & eh_1 ^ abc_0 & eg_1 ^ abc_0 & efh_1 ^ abc_0 & efg_1 ^ abc_0 & efgh_1 ^ abcd_0 & h_1 ^ abcd_0 & f_1 ^ abcd_0 & fg_1 ^ abcd_0 & e_1 ^ abcd_0 & egh_1 ^ abcd_0 & ef_1 ^ abcd_0 & efh_1 ;
        assign f3_10 = d_1 & gh_0 ^ d_1 & fh_0 ^ d_1 & fgh_0 ^ d_1 & eh_0 ^ d_1 & eg_0 ^ d_1 & ef_0 ^ d_1 & efgh_0 ^ c_1 & gh_0 ^ c_1 & fg_0 ^ c_1 & fgh_0 ^ c_1 & ef_0 ^ c_1 & efg_0 ^ c_1 & efgh_0 ^ cd_1 & h_0 ^ cd_1 & f_0 ^ cd_1 & fg_0 ^ cd_1 & eg_0 ^ cd_1 & egh_0 ^ cd_1 & ef_0 ^ cd_1 & efh_0 ^ b_1 & gh_0 ^ b_1 & fh_0 ^ b_1 & fg_0 ^ b_1 & e_0 ^ b_1 & eh_0 ^ b_1 & egh_0 ^ b_1 & efg_0 ^ bd_1 & h_0 ^ bd_1 & gh_0 ^ bd_1 & fh_0 ^ bd_1 & eh_0 ^ bd_1 & eg_0 ^ bd_1 & egh_0 ^ bd_1 & efgh_0 ^ bc_1 & g_0 ^ bc_1 & gh_0 ^ bc_1 & fh_0 ^ bc_1 & fgh_0 ^ bc_1 & e_0 ^ bc_1 & eg_0 ^ bc_1 & egh_0 ^ bc_1 & efh_0 ^ bc_1 & efg_0 ^ bc_1 & efgh_0 ^ bcd_1 & h_0 ^ bcd_1 & g_0 ^ bcd_1 & f_0 ^ bcd_1 & fh_0 ^ bcd_1 & fg_0 ^ bcd_1 & e_0 ^ bcd_1 & eh_0 ^ bcd_1 & ef_0 ^ bcd_1 & efg_0 ^ bcd_1 & efgh_0 ^ a_1 & h_0 ^ a_1 & g_0 ^ a_1 & gh_0 ^ a_1 & fh_0 ^ a_1 & fg_0 ^ a_1 & e_0 ^ a_1 & eh_0 ^ a_1 & ef_0 ^ a_1 & efh_0 ^ a_1 & efg_0 ^ a_1 & efgh_0 ^ ad_1 & fh_0 ^ ad_1 & fg_0 ^ ad_1 & fgh_0 ^ ad_1 & e_0 ^ ad_1 & eg_0 ^ ad_1 & egh_0 ^ ad_1 & efgh_0 ^ ac_1 & f_0 ^ ac_1 & fg_0 ^ ac_1 & fgh_0 ^ ac_1 & e_0 ^ ac_1 & efh_0 ^ ac_1 & efgh_0 ^ acd_1 & g_0 ^ acd_1 & gh_0 ^ acd_1 & f_0 ^ acd_1 & fh_0 ^ acd_1 & fgh_0 ^ acd_1 & eh_0 ^ acd_1 & egh_0 ^ acd_1 & ef_0 ^ acd_1 & efg_0 ^ ab_1 & gh_0 ^ ab_1 & fh_0 ^ ab_1 & fg_0 ^ ab_1 & eh_0 ^ ab_1 & efh_0 ^ ab_1 & efgh_0 ^ abd_1 & g_0 ^ abd_1 & f_0 ^ abd_1 & fgh_0 ^ abd_1 & e_0 ^ abd_1 & eh_0 ^ abd_1 & eg_0 ^ abd_1 & efh_0 ^ abd_1 & efg_0 ^ abc_1 & h_0 ^ abc_1 & g_0 ^ abc_1 & gh_0 ^ abc_1 & fh_0 ^ abc_1 & fg_0 ^ abc_1 & e_0 ^ abc_1 & eh_0 ^ abc_1 & eg_0 ^ abc_1 & efh_0 ^ abc_1 & efg_0 ^ abc_1 & efgh_0 ^ abcd_1 & h_0 ^ abcd_1 & f_0 ^ abcd_1 & fg_0 ^ abcd_1 & e_0 ^ abcd_1 & egh_0 ^ abcd_1 & ef_0 ^ abcd_1 & efh_0 ;
        assign f3_11 = h_1 ^ fg_1 ^ eh_1 ^ egh_1 ^ ef_1 ^ efh_1 ^ efg_1 ^ efgh_1 ^ d_1 ^ d_1 & gh_1 ^ d_1 & fh_1 ^ d_1 & fgh_1 ^ d_1 & eh_1 ^ d_1 & eg_1 ^ d_1 & ef_1 ^ d_1 & efgh_1 ^ c_1 & gh_1 ^ c_1 & fg_1 ^ c_1 & fgh_1 ^ c_1 & ef_1 ^ c_1 & efg_1 ^ c_1 & efgh_1 ^ cd_1 ^ cd_1 & h_1 ^ cd_1 & f_1 ^ cd_1 & fg_1 ^ cd_1 & eg_1 ^ cd_1 & egh_1 ^ cd_1 & ef_1 ^ cd_1 & efh_1 ^ b_1 ^ b_1 & gh_1 ^ b_1 & fh_1 ^ b_1 & fg_1 ^ b_1 & e_1 ^ b_1 & eh_1 ^ b_1 & egh_1 ^ b_1 & efg_1 ^ bd_1 & h_1 ^ bd_1 & gh_1 ^ bd_1 & fh_1 ^ bd_1 & eh_1 ^ bd_1 & eg_1 ^ bd_1 & egh_1 ^ bd_1 & efgh_1 ^ bc_1 ^ bc_1 & g_1 ^ bc_1 & gh_1 ^ bc_1 & fh_1 ^ bc_1 & fgh_1 ^ bc_1 & e_1 ^ bc_1 & eg_1 ^ bc_1 & egh_1 ^ bc_1 & efh_1 ^ bc_1 & efg_1 ^ bc_1 & efgh_1 ^ bcd_1 & h_1 ^ bcd_1 & g_1 ^ bcd_1 & f_1 ^ bcd_1 & fh_1 ^ bcd_1 & fg_1 ^ bcd_1 & e_1 ^ bcd_1 & eh_1 ^ bcd_1 & ef_1 ^ bcd_1 & efg_1 ^ bcd_1 & efgh_1 ^ a_1 ^ a_1 & h_1 ^ a_1 & g_1 ^ a_1 & gh_1 ^ a_1 & fh_1 ^ a_1 & fg_1 ^ a_1 & e_1 ^ a_1 & eh_1 ^ a_1 & ef_1 ^ a_1 & efh_1 ^ a_1 & efg_1 ^ a_1 & efgh_1 ^ ad_1 & fh_1 ^ ad_1 & fg_1 ^ ad_1 & fgh_1 ^ ad_1 & e_1 ^ ad_1 & eg_1 ^ ad_1 & egh_1 ^ ad_1 & efgh_1 ^ ac_1 ^ ac_1 & f_1 ^ ac_1 & fg_1 ^ ac_1 & fgh_1 ^ ac_1 & e_1 ^ ac_1 & efh_1 ^ ac_1 & efgh_1 ^ acd_1 & g_1 ^ acd_1 & gh_1 ^ acd_1 & f_1 ^ acd_1 & fh_1 ^ acd_1 & fgh_1 ^ acd_1 & eh_1 ^ acd_1 & egh_1 ^ acd_1 & ef_1 ^ acd_1 & efg_1 ^ ab_1 ^ ab_1 & gh_1 ^ ab_1 & fh_1 ^ ab_1 & fg_1 ^ ab_1 & eh_1 ^ ab_1 & efh_1 ^ ab_1 & efgh_1 ^ abd_1 & g_1 ^ abd_1 & f_1 ^ abd_1 & fgh_1 ^ abd_1 & e_1 ^ abd_1 & eh_1 ^ abd_1 & eg_1 ^ abd_1 & efh_1 ^ abd_1 & efg_1 ^ abc_1 ^ abc_1 & h_1 ^ abc_1 & g_1 ^ abc_1 & gh_1 ^ abc_1 & fh_1 ^ abc_1 & fg_1 ^ abc_1 & e_1 ^ abc_1 & eh_1 ^ abc_1 & eg_1 ^ abc_1 & efh_1 ^ abc_1 & efg_1 ^ abc_1 & efgh_1 ^ abcd_1 ^ abcd_1 & h_1 ^ abcd_1 & f_1 ^ abcd_1 & fg_1 ^ abcd_1 & e_1 ^ abcd_1 & egh_1 ^ abcd_1 & ef_1 ^ abcd_1 & efh_1 ;
        wire f3_00_reg;
        Register # (1) inst_inner_f3_00 (f3_00, clk, f3_00_reg);
        wire f3_01_reg;
        Register # (1) inst_cross_f3_01 (f3_01 ^ r_cross[3], clk, f3_01_reg);
        wire f3_10_reg;
        Register # (1) inst_cross_f3_10 (f3_10 ^ r_cross[3], clk, f3_10_reg);
        wire f3_11_reg;
        Register # (1) inst_inner_f3_11 (f3_11, clk, f3_11_reg);
        //////////////
        
        assign f4_00 = h_0 ^ g_0 ^ gh_0 ^ f_0 ^ e_0 ^ ef_0 ^ efh_0 ^ d_0 & h_0 ^ d_0 & g_0 ^ d_0 & fg_0 ^ d_0 & e_0 ^ d_0 & eh_0 ^ d_0 & ef_0 ^ d_0 & efh_0 ^ d_0 & efg_0 ^ d_0 & efgh_0 ^ c_0 ^ c_0 & h_0 ^ c_0 & g_0 ^ c_0 & f_0 ^ c_0 & e_0 ^ c_0 & eh_0 ^ c_0 & eg_0 ^ c_0 & egh_0 ^ c_0 & ef_0 ^ c_0 & efg_0 ^ cd_0 ^ cd_0 & h_0 ^ cd_0 & g_0 ^ cd_0 & gh_0 ^ cd_0 & f_0 ^ cd_0 & fgh_0 ^ cd_0 & e_0 ^ cd_0 & eh_0 ^ cd_0 & eg_0 ^ cd_0 & efh_0 ^ cd_0 & efgh_0 ^ b_0 & h_0 ^ b_0 & g_0 ^ b_0 & fh_0 ^ b_0 & fgh_0 ^ b_0 & egh_0 ^ b_0 & ef_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & h_0 ^ bd_0 & gh_0 ^ bd_0 & fg_0 ^ bd_0 & e_0 ^ bd_0 & eh_0 ^ bd_0 & egh_0 ^ bd_0 & efh_0 ^ bd_0 & efg_0 ^ bc_0 & gh_0 ^ bc_0 & f_0 ^ bc_0 & e_0 ^ bc_0 & eh_0 ^ bc_0 & ef_0 ^ bc_0 & efh_0 ^ bc_0 & efg_0 ^ bc_0 & efgh_0 ^ bcd_0 & h_0 ^ bcd_0 & gh_0 ^ bcd_0 & fg_0 ^ bcd_0 & fgh_0 ^ bcd_0 & eg_0 ^ bcd_0 & egh_0 ^ bcd_0 & ef_0 ^ bcd_0 & efg_0 ^ a_0 & h_0 ^ a_0 & e_0 ^ a_0 & egh_0 ^ a_0 & efgh_0 ^ ad_0 & h_0 ^ ad_0 & f_0 ^ ad_0 & e_0 ^ ad_0 & eh_0 ^ ad_0 & eg_0 ^ ad_0 & ef_0 ^ ad_0 & efgh_0 ^ ac_0 ^ ac_0 & g_0 ^ ac_0 & gh_0 ^ ac_0 & fh_0 ^ ac_0 & fg_0 ^ ac_0 & fgh_0 ^ ac_0 & e_0 ^ ac_0 & eh_0 ^ ac_0 & egh_0 ^ ac_0 & ef_0 ^ ac_0 & efh_0 ^ ac_0 & efg_0 ^ acd_0 ^ acd_0 & fg_0 ^ acd_0 & e_0 ^ acd_0 & eg_0 ^ acd_0 & ef_0 ^ acd_0 & efh_0 ^ acd_0 & efg_0 ^ acd_0 & efgh_0 ^ ab_0 ^ ab_0 & h_0 ^ ab_0 & g_0 ^ ab_0 & gh_0 ^ ab_0 & f_0 ^ ab_0 & fg_0 ^ ab_0 & fgh_0 ^ ab_0 & e_0 ^ ab_0 & eh_0 ^ ab_0 & egh_0 ^ abd_0 ^ abd_0 & h_0 ^ abd_0 & fh_0 ^ abd_0 & e_0 ^ abd_0 & eh_0 ^ abd_0 & ef_0 ^ abd_0 & efg_0 ^ abd_0 & efgh_0 ^ abc_0 ^ abc_0 & gh_0 ^ abc_0 & fg_0 ^ abc_0 & e_0 ^ abc_0 & eh_0 ^ abc_0 & eg_0 ^ abc_0 & efg_0 ^ abcd_0 & h_0 ^ abcd_0 & g_0 ^ abcd_0 & f_0 ^ abcd_0 & e_0 ^ abcd_0 & eh_0 ^ abcd_0 & efh_0 ;
        assign f4_01 = d_0 & h_1 ^ d_0 & g_1 ^ d_0 & fg_1 ^ d_0 & e_1 ^ d_0 & eh_1 ^ d_0 & ef_1 ^ d_0 & efh_1 ^ d_0 & efg_1 ^ d_0 & efgh_1 ^ c_0 & h_1 ^ c_0 & g_1 ^ c_0 & f_1 ^ c_0 & e_1 ^ c_0 & eh_1 ^ c_0 & eg_1 ^ c_0 & egh_1 ^ c_0 & ef_1 ^ c_0 & efg_1 ^ cd_0 & h_1 ^ cd_0 & g_1 ^ cd_0 & gh_1 ^ cd_0 & f_1 ^ cd_0 & fgh_1 ^ cd_0 & e_1 ^ cd_0 & eh_1 ^ cd_0 & eg_1 ^ cd_0 & efh_1 ^ cd_0 & efgh_1 ^ b_0 & h_1 ^ b_0 & g_1 ^ b_0 & fh_1 ^ b_0 & fgh_1 ^ b_0 & egh_1 ^ b_0 & ef_1 ^ b_0 & efgh_1 ^ bd_0 & h_1 ^ bd_0 & gh_1 ^ bd_0 & fg_1 ^ bd_0 & e_1 ^ bd_0 & eh_1 ^ bd_0 & egh_1 ^ bd_0 & efh_1 ^ bd_0 & efg_1 ^ bc_0 & gh_1 ^ bc_0 & f_1 ^ bc_0 & e_1 ^ bc_0 & eh_1 ^ bc_0 & ef_1 ^ bc_0 & efh_1 ^ bc_0 & efg_1 ^ bc_0 & efgh_1 ^ bcd_0 & h_1 ^ bcd_0 & gh_1 ^ bcd_0 & fg_1 ^ bcd_0 & fgh_1 ^ bcd_0 & eg_1 ^ bcd_0 & egh_1 ^ bcd_0 & ef_1 ^ bcd_0 & efg_1 ^ a_0 & h_1 ^ a_0 & e_1 ^ a_0 & egh_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & f_1 ^ ad_0 & e_1 ^ ad_0 & eh_1 ^ ad_0 & eg_1 ^ ad_0 & ef_1 ^ ad_0 & efgh_1 ^ ac_0 & g_1 ^ ac_0 & gh_1 ^ ac_0 & fh_1 ^ ac_0 & fg_1 ^ ac_0 & fgh_1 ^ ac_0 & e_1 ^ ac_0 & eh_1 ^ ac_0 & egh_1 ^ ac_0 & ef_1 ^ ac_0 & efh_1 ^ ac_0 & efg_1 ^ acd_0 & fg_1 ^ acd_0 & e_1 ^ acd_0 & eg_1 ^ acd_0 & ef_1 ^ acd_0 & efh_1 ^ acd_0 & efg_1 ^ acd_0 & efgh_1 ^ ab_0 & h_1 ^ ab_0 & g_1 ^ ab_0 & gh_1 ^ ab_0 & f_1 ^ ab_0 & fg_1 ^ ab_0 & fgh_1 ^ ab_0 & e_1 ^ ab_0 & eh_1 ^ ab_0 & egh_1 ^ abd_0 & h_1 ^ abd_0 & fh_1 ^ abd_0 & e_1 ^ abd_0 & eh_1 ^ abd_0 & ef_1 ^ abd_0 & efg_1 ^ abd_0 & efgh_1 ^ abc_0 & gh_1 ^ abc_0 & fg_1 ^ abc_0 & e_1 ^ abc_0 & eh_1 ^ abc_0 & eg_1 ^ abc_0 & efg_1 ^ abcd_0 & h_1 ^ abcd_0 & g_1 ^ abcd_0 & f_1 ^ abcd_0 & e_1 ^ abcd_0 & eh_1 ^ abcd_0 & efh_1 ;
        assign f4_10 = d_1 & h_0 ^ d_1 & g_0 ^ d_1 & fg_0 ^ d_1 & e_0 ^ d_1 & eh_0 ^ d_1 & ef_0 ^ d_1 & efh_0 ^ d_1 & efg_0 ^ d_1 & efgh_0 ^ c_1 & h_0 ^ c_1 & g_0 ^ c_1 & f_0 ^ c_1 & e_0 ^ c_1 & eh_0 ^ c_1 & eg_0 ^ c_1 & egh_0 ^ c_1 & ef_0 ^ c_1 & efg_0 ^ cd_1 & h_0 ^ cd_1 & g_0 ^ cd_1 & gh_0 ^ cd_1 & f_0 ^ cd_1 & fgh_0 ^ cd_1 & e_0 ^ cd_1 & eh_0 ^ cd_1 & eg_0 ^ cd_1 & efh_0 ^ cd_1 & efgh_0 ^ b_1 & h_0 ^ b_1 & g_0 ^ b_1 & fh_0 ^ b_1 & fgh_0 ^ b_1 & egh_0 ^ b_1 & ef_0 ^ b_1 & efgh_0 ^ bd_1 & h_0 ^ bd_1 & gh_0 ^ bd_1 & fg_0 ^ bd_1 & e_0 ^ bd_1 & eh_0 ^ bd_1 & egh_0 ^ bd_1 & efh_0 ^ bd_1 & efg_0 ^ bc_1 & gh_0 ^ bc_1 & f_0 ^ bc_1 & e_0 ^ bc_1 & eh_0 ^ bc_1 & ef_0 ^ bc_1 & efh_0 ^ bc_1 & efg_0 ^ bc_1 & efgh_0 ^ bcd_1 & h_0 ^ bcd_1 & gh_0 ^ bcd_1 & fg_0 ^ bcd_1 & fgh_0 ^ bcd_1 & eg_0 ^ bcd_1 & egh_0 ^ bcd_1 & ef_0 ^ bcd_1 & efg_0 ^ a_1 & h_0 ^ a_1 & e_0 ^ a_1 & egh_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & f_0 ^ ad_1 & e_0 ^ ad_1 & eh_0 ^ ad_1 & eg_0 ^ ad_1 & ef_0 ^ ad_1 & efgh_0 ^ ac_1 & g_0 ^ ac_1 & gh_0 ^ ac_1 & fh_0 ^ ac_1 & fg_0 ^ ac_1 & fgh_0 ^ ac_1 & e_0 ^ ac_1 & eh_0 ^ ac_1 & egh_0 ^ ac_1 & ef_0 ^ ac_1 & efh_0 ^ ac_1 & efg_0 ^ acd_1 & fg_0 ^ acd_1 & e_0 ^ acd_1 & eg_0 ^ acd_1 & ef_0 ^ acd_1 & efh_0 ^ acd_1 & efg_0 ^ acd_1 & efgh_0 ^ ab_1 & h_0 ^ ab_1 & g_0 ^ ab_1 & gh_0 ^ ab_1 & f_0 ^ ab_1 & fg_0 ^ ab_1 & fgh_0 ^ ab_1 & e_0 ^ ab_1 & eh_0 ^ ab_1 & egh_0 ^ abd_1 & h_0 ^ abd_1 & fh_0 ^ abd_1 & e_0 ^ abd_1 & eh_0 ^ abd_1 & ef_0 ^ abd_1 & efg_0 ^ abd_1 & efgh_0 ^ abc_1 & gh_0 ^ abc_1 & fg_0 ^ abc_1 & e_0 ^ abc_1 & eh_0 ^ abc_1 & eg_0 ^ abc_1 & efg_0 ^ abcd_1 & h_0 ^ abcd_1 & g_0 ^ abcd_1 & f_0 ^ abcd_1 & e_0 ^ abcd_1 & eh_0 ^ abcd_1 & efh_0 ;
        assign f4_11 = h_1 ^ g_1 ^ gh_1 ^ f_1 ^ e_1 ^ ef_1 ^ efh_1 ^ d_1 & h_1 ^ d_1 & g_1 ^ d_1 & fg_1 ^ d_1 & e_1 ^ d_1 & eh_1 ^ d_1 & ef_1 ^ d_1 & efh_1 ^ d_1 & efg_1 ^ d_1 & efgh_1 ^ c_1 ^ c_1 & h_1 ^ c_1 & g_1 ^ c_1 & f_1 ^ c_1 & e_1 ^ c_1 & eh_1 ^ c_1 & eg_1 ^ c_1 & egh_1 ^ c_1 & ef_1 ^ c_1 & efg_1 ^ cd_1 ^ cd_1 & h_1 ^ cd_1 & g_1 ^ cd_1 & gh_1 ^ cd_1 & f_1 ^ cd_1 & fgh_1 ^ cd_1 & e_1 ^ cd_1 & eh_1 ^ cd_1 & eg_1 ^ cd_1 & efh_1 ^ cd_1 & efgh_1 ^ b_1 & h_1 ^ b_1 & g_1 ^ b_1 & fh_1 ^ b_1 & fgh_1 ^ b_1 & egh_1 ^ b_1 & ef_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & h_1 ^ bd_1 & gh_1 ^ bd_1 & fg_1 ^ bd_1 & e_1 ^ bd_1 & eh_1 ^ bd_1 & egh_1 ^ bd_1 & efh_1 ^ bd_1 & efg_1 ^ bc_1 & gh_1 ^ bc_1 & f_1 ^ bc_1 & e_1 ^ bc_1 & eh_1 ^ bc_1 & ef_1 ^ bc_1 & efh_1 ^ bc_1 & efg_1 ^ bc_1 & efgh_1 ^ bcd_1 & h_1 ^ bcd_1 & gh_1 ^ bcd_1 & fg_1 ^ bcd_1 & fgh_1 ^ bcd_1 & eg_1 ^ bcd_1 & egh_1 ^ bcd_1 & ef_1 ^ bcd_1 & efg_1 ^ a_1 & h_1 ^ a_1 & e_1 ^ a_1 & egh_1 ^ a_1 & efgh_1 ^ ad_1 & h_1 ^ ad_1 & f_1 ^ ad_1 & e_1 ^ ad_1 & eh_1 ^ ad_1 & eg_1 ^ ad_1 & ef_1 ^ ad_1 & efgh_1 ^ ac_1 ^ ac_1 & g_1 ^ ac_1 & gh_1 ^ ac_1 & fh_1 ^ ac_1 & fg_1 ^ ac_1 & fgh_1 ^ ac_1 & e_1 ^ ac_1 & eh_1 ^ ac_1 & egh_1 ^ ac_1 & ef_1 ^ ac_1 & efh_1 ^ ac_1 & efg_1 ^ acd_1 ^ acd_1 & fg_1 ^ acd_1 & e_1 ^ acd_1 & eg_1 ^ acd_1 & ef_1 ^ acd_1 & efh_1 ^ acd_1 & efg_1 ^ acd_1 & efgh_1 ^ ab_1 ^ ab_1 & h_1 ^ ab_1 & g_1 ^ ab_1 & gh_1 ^ ab_1 & f_1 ^ ab_1 & fg_1 ^ ab_1 & fgh_1 ^ ab_1 & e_1 ^ ab_1 & eh_1 ^ ab_1 & egh_1 ^ abd_1 ^ abd_1 & h_1 ^ abd_1 & fh_1 ^ abd_1 & e_1 ^ abd_1 & eh_1 ^ abd_1 & ef_1 ^ abd_1 & efg_1 ^ abd_1 & efgh_1 ^ abc_1 ^ abc_1 & gh_1 ^ abc_1 & fg_1 ^ abc_1 & e_1 ^ abc_1 & eh_1 ^ abc_1 & eg_1 ^ abc_1 & efg_1 ^ abcd_1 & h_1 ^ abcd_1 & g_1 ^ abcd_1 & f_1 ^ abcd_1 & e_1 ^ abcd_1 & eh_1 ^ abcd_1 & efh_1 ;
        wire f4_00_reg;
        Register # (1) inst_inner_f4_00 (f4_00, clk, f4_00_reg);
        wire f4_01_reg;
        Register # (1) inst_cross_f4_01 (f4_01 ^ r_cross[4], clk, f4_01_reg);
        wire f4_10_reg;
        Register # (1) inst_cross_f4_10 (f4_10 ^ r_cross[4], clk, f4_10_reg);
        wire f4_11_reg;
        Register # (1) inst_inner_f4_11 (f4_11, clk, f4_11_reg);
        /////////////
        
        assign f5_00 = fgh_0 ^ eh_0 ^ egh_0 ^ efgh_0 ^ d_0 ^ d_0 & gh_0 ^ d_0 & f_0 ^ d_0 & fh_0 ^ d_0 & fg_0 ^ d_0 & e_0 ^ d_0 & egh_0 ^ d_0 & efh_0 ^ d_0 & efgh_0 ^ c_0 & g_0 ^ c_0 & gh_0 ^ c_0 & fg_0 ^ c_0 & fgh_0 ^ c_0 & eh_0 ^ c_0 & eg_0 ^ c_0 & efh_0 ^ c_0 & efg_0 ^ c_0 & efgh_0 ^ cd_0 & gh_0 ^ cd_0 & f_0 ^ cd_0 & fh_0 ^ cd_0 & fg_0 ^ cd_0 & fgh_0 ^ cd_0 & e_0 ^ cd_0 & ef_0 ^ cd_0 & efgh_0 ^ b_0 ^ b_0 & g_0 ^ b_0 & gh_0 ^ b_0 & fh_0 ^ b_0 & fg_0 ^ b_0 & eg_0 ^ b_0 & ef_0 ^ b_0 & efg_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & g_0 ^ bd_0 & gh_0 ^ bd_0 & fgh_0 ^ bd_0 & eg_0 ^ bd_0 & ef_0 ^ bd_0 & efg_0 ^ bc_0 & h_0 ^ bc_0 & g_0 ^ bc_0 & gh_0 ^ bc_0 & eg_0 ^ bc_0 & ef_0 ^ bc_0 & efgh_0 ^ bcd_0 & gh_0 ^ bcd_0 & fg_0 ^ bcd_0 & fgh_0 ^ bcd_0 & e_0 ^ bcd_0 & eh_0 ^ bcd_0 & eg_0 ^ bcd_0 & ef_0 ^ a_0 ^ a_0 & gh_0 ^ a_0 & eg_0 ^ a_0 & egh_0 ^ a_0 & ef_0 ^ a_0 & efgh_0 ^ ad_0 & h_0 ^ ad_0 & g_0 ^ ad_0 & gh_0 ^ ad_0 & f_0 ^ ad_0 & fg_0 ^ ad_0 & eh_0 ^ ad_0 & eg_0 ^ ad_0 & ef_0 ^ ad_0 & efh_0 ^ ad_0 & efg_0 ^ ac_0 ^ ac_0 & g_0 ^ ac_0 & gh_0 ^ ac_0 & f_0 ^ ac_0 & e_0 ^ ac_0 & eg_0 ^ ac_0 & egh_0 ^ ac_0 & efh_0 ^ ac_0 & efgh_0 ^ acd_0 ^ acd_0 & g_0 ^ acd_0 & gh_0 ^ acd_0 & f_0 ^ acd_0 & fh_0 ^ acd_0 & fgh_0 ^ acd_0 & e_0 ^ acd_0 & eh_0 ^ ab_0 & g_0 ^ ab_0 & f_0 ^ ab_0 & fgh_0 ^ ab_0 & efh_0 ^ abd_0 & h_0 ^ abd_0 & gh_0 ^ abd_0 & e_0 ^ abd_0 & eg_0 ^ abd_0 & efh_0 ^ abd_0 & efg_0 ^ abc_0 ^ abc_0 & h_0 ^ abc_0 & gh_0 ^ abc_0 & ef_0 ^ abc_0 & efg_0 ^ abc_0 & efgh_0 ^ abcd_0 & h_0 ^ abcd_0 & f_0 ^ abcd_0 & fh_0 ^ abcd_0 & fg_0 ^ abcd_0 & fgh_0 ;
        assign f5_01 = d_0 & gh_1 ^ d_0 & f_1 ^ d_0 & fh_1 ^ d_0 & fg_1 ^ d_0 & e_1 ^ d_0 & egh_1 ^ d_0 & efh_1 ^ d_0 & efgh_1 ^ c_0 & g_1 ^ c_0 & gh_1 ^ c_0 & fg_1 ^ c_0 & fgh_1 ^ c_0 & eh_1 ^ c_0 & eg_1 ^ c_0 & efh_1 ^ c_0 & efg_1 ^ c_0 & efgh_1 ^ cd_0 & gh_1 ^ cd_0 & f_1 ^ cd_0 & fh_1 ^ cd_0 & fg_1 ^ cd_0 & fgh_1 ^ cd_0 & e_1 ^ cd_0 & ef_1 ^ cd_0 & efgh_1 ^ b_0 & g_1 ^ b_0 & gh_1 ^ b_0 & fh_1 ^ b_0 & fg_1 ^ b_0 & eg_1 ^ b_0 & ef_1 ^ b_0 & efg_1 ^ b_0 & efgh_1 ^ bd_0 & g_1 ^ bd_0 & gh_1 ^ bd_0 & fgh_1 ^ bd_0 & eg_1 ^ bd_0 & ef_1 ^ bd_0 & efg_1 ^ bc_0 & h_1 ^ bc_0 & g_1 ^ bc_0 & gh_1 ^ bc_0 & eg_1 ^ bc_0 & ef_1 ^ bc_0 & efgh_1 ^ bcd_0 & gh_1 ^ bcd_0 & fg_1 ^ bcd_0 & fgh_1 ^ bcd_0 & e_1 ^ bcd_0 & eh_1 ^ bcd_0 & eg_1 ^ bcd_0 & ef_1 ^ a_0 & gh_1 ^ a_0 & eg_1 ^ a_0 & egh_1 ^ a_0 & ef_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & g_1 ^ ad_0 & gh_1 ^ ad_0 & f_1 ^ ad_0 & fg_1 ^ ad_0 & eh_1 ^ ad_0 & eg_1 ^ ad_0 & ef_1 ^ ad_0 & efh_1 ^ ad_0 & efg_1 ^ ac_0 & g_1 ^ ac_0 & gh_1 ^ ac_0 & f_1 ^ ac_0 & e_1 ^ ac_0 & eg_1 ^ ac_0 & egh_1 ^ ac_0 & efh_1 ^ ac_0 & efgh_1 ^ acd_0 & g_1 ^ acd_0 & gh_1 ^ acd_0 & f_1 ^ acd_0 & fh_1 ^ acd_0 & fgh_1 ^ acd_0 & e_1 ^ acd_0 & eh_1 ^ ab_0 & g_1 ^ ab_0 & f_1 ^ ab_0 & fgh_1 ^ ab_0 & efh_1 ^ abd_0 & h_1 ^ abd_0 & gh_1 ^ abd_0 & e_1 ^ abd_0 & eg_1 ^ abd_0 & efh_1 ^ abd_0 & efg_1 ^ abc_0 & h_1 ^ abc_0 & gh_1 ^ abc_0 & ef_1 ^ abc_0 & efg_1 ^ abc_0 & efgh_1 ^ abcd_0 & h_1 ^ abcd_0 & f_1 ^ abcd_0 & fh_1 ^ abcd_0 & fg_1 ^ abcd_0 & fgh_1 ;
        assign f5_10 = d_1 & gh_0 ^ d_1 & f_0 ^ d_1 & fh_0 ^ d_1 & fg_0 ^ d_1 & e_0 ^ d_1 & egh_0 ^ d_1 & efh_0 ^ d_1 & efgh_0 ^ c_1 & g_0 ^ c_1 & gh_0 ^ c_1 & fg_0 ^ c_1 & fgh_0 ^ c_1 & eh_0 ^ c_1 & eg_0 ^ c_1 & efh_0 ^ c_1 & efg_0 ^ c_1 & efgh_0 ^ cd_1 & gh_0 ^ cd_1 & f_0 ^ cd_1 & fh_0 ^ cd_1 & fg_0 ^ cd_1 & fgh_0 ^ cd_1 & e_0 ^ cd_1 & ef_0 ^ cd_1 & efgh_0 ^ b_1 & g_0 ^ b_1 & gh_0 ^ b_1 & fh_0 ^ b_1 & fg_0 ^ b_1 & eg_0 ^ b_1 & ef_0 ^ b_1 & efg_0 ^ b_1 & efgh_0 ^ bd_1 & g_0 ^ bd_1 & gh_0 ^ bd_1 & fgh_0 ^ bd_1 & eg_0 ^ bd_1 & ef_0 ^ bd_1 & efg_0 ^ bc_1 & h_0 ^ bc_1 & g_0 ^ bc_1 & gh_0 ^ bc_1 & eg_0 ^ bc_1 & ef_0 ^ bc_1 & efgh_0 ^ bcd_1 & gh_0 ^ bcd_1 & fg_0 ^ bcd_1 & fgh_0 ^ bcd_1 & e_0 ^ bcd_1 & eh_0 ^ bcd_1 & eg_0 ^ bcd_1 & ef_0 ^ a_1 & gh_0 ^ a_1 & eg_0 ^ a_1 & egh_0 ^ a_1 & ef_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & g_0 ^ ad_1 & gh_0 ^ ad_1 & f_0 ^ ad_1 & fg_0 ^ ad_1 & eh_0 ^ ad_1 & eg_0 ^ ad_1 & ef_0 ^ ad_1 & efh_0 ^ ad_1 & efg_0 ^ ac_1 & g_0 ^ ac_1 & gh_0 ^ ac_1 & f_0 ^ ac_1 & e_0 ^ ac_1 & eg_0 ^ ac_1 & egh_0 ^ ac_1 & efh_0 ^ ac_1 & efgh_0 ^ acd_1 & g_0 ^ acd_1 & gh_0 ^ acd_1 & f_0 ^ acd_1 & fh_0 ^ acd_1 & fgh_0 ^ acd_1 & e_0 ^ acd_1 & eh_0 ^ ab_1 & g_0 ^ ab_1 & f_0 ^ ab_1 & fgh_0 ^ ab_1 & efh_0 ^ abd_1 & h_0 ^ abd_1 & gh_0 ^ abd_1 & e_0 ^ abd_1 & eg_0 ^ abd_1 & efh_0 ^ abd_1 & efg_0 ^ abc_1 & h_0 ^ abc_1 & gh_0 ^ abc_1 & ef_0 ^ abc_1 & efg_0 ^ abc_1 & efgh_0 ^ abcd_1 & h_0 ^ abcd_1 & f_0 ^ abcd_1 & fh_0 ^ abcd_1 & fg_0 ^ abcd_1 & fgh_0 ;
        assign f5_11 = fgh_1 ^ eh_1 ^ egh_1 ^ efgh_1 ^ d_1 ^ d_1 & gh_1 ^ d_1 & f_1 ^ d_1 & fh_1 ^ d_1 & fg_1 ^ d_1 & e_1 ^ d_1 & egh_1 ^ d_1 & efh_1 ^ d_1 & efgh_1 ^ c_1 & g_1 ^ c_1 & gh_1 ^ c_1 & fg_1 ^ c_1 & fgh_1 ^ c_1 & eh_1 ^ c_1 & eg_1 ^ c_1 & efh_1 ^ c_1 & efg_1 ^ c_1 & efgh_1 ^ cd_1 & gh_1 ^ cd_1 & f_1 ^ cd_1 & fh_1 ^ cd_1 & fg_1 ^ cd_1 & fgh_1 ^ cd_1 & e_1 ^ cd_1 & ef_1 ^ cd_1 & efgh_1 ^ b_1 ^ b_1 & g_1 ^ b_1 & gh_1 ^ b_1 & fh_1 ^ b_1 & fg_1 ^ b_1 & eg_1 ^ b_1 & ef_1 ^ b_1 & efg_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & g_1 ^ bd_1 & gh_1 ^ bd_1 & fgh_1 ^ bd_1 & eg_1 ^ bd_1 & ef_1 ^ bd_1 & efg_1 ^ bc_1 & h_1 ^ bc_1 & g_1 ^ bc_1 & gh_1 ^ bc_1 & eg_1 ^ bc_1 & ef_1 ^ bc_1 & efgh_1 ^ bcd_1 & gh_1 ^ bcd_1 & fg_1 ^ bcd_1 & fgh_1 ^ bcd_1 & e_1 ^ bcd_1 & eh_1 ^ bcd_1 & eg_1 ^ bcd_1 & ef_1 ^ a_1 ^ a_1 & gh_1 ^ a_1 & eg_1 ^ a_1 & egh_1 ^ a_1 & ef_1 ^ a_1 & efgh_1 ^ ad_1 & h_1 ^ ad_1 & g_1 ^ ad_1 & gh_1 ^ ad_1 & f_1 ^ ad_1 & fg_1 ^ ad_1 & eh_1 ^ ad_1 & eg_1 ^ ad_1 & ef_1 ^ ad_1 & efh_1 ^ ad_1 & efg_1 ^ ac_1 ^ ac_1 & g_1 ^ ac_1 & gh_1 ^ ac_1 & f_1 ^ ac_1 & e_1 ^ ac_1 & eg_1 ^ ac_1 & egh_1 ^ ac_1 & efh_1 ^ ac_1 & efgh_1 ^ acd_1 ^ acd_1 & g_1 ^ acd_1 & gh_1 ^ acd_1 & f_1 ^ acd_1 & fh_1 ^ acd_1 & fgh_1 ^ acd_1 & e_1 ^ acd_1 & eh_1 ^ ab_1 & g_1 ^ ab_1 & f_1 ^ ab_1 & fgh_1 ^ ab_1 & efh_1 ^ abd_1 & h_1 ^ abd_1 & gh_1 ^ abd_1 & e_1 ^ abd_1 & eg_1 ^ abd_1 & efh_1 ^ abd_1 & efg_1 ^ abc_1 ^ abc_1 & h_1 ^ abc_1 & gh_1 ^ abc_1 & ef_1 ^ abc_1 & efg_1 ^ abc_1 & efgh_1 ^ abcd_1 & h_1 ^ abcd_1 & f_1 ^ abcd_1 & fh_1 ^ abcd_1 & fg_1 ^ abcd_1 & fgh_1 ;
        wire f5_00_reg;
        Register # (1) inst_inner_f5_00 (f5_00, clk, f5_00_reg);
        wire f5_01_reg;
        Register # (1) inst_cross_f5_01 (f5_01 ^ r_cross[5], clk, f5_01_reg);
        wire f5_10_reg;
        Register # (1) inst_cross_f5_10 (f5_10 ^ r_cross[5], clk, f5_10_reg);
        wire f5_11_reg;
        Register # (1) inst_inner_f5_11 (f5_11, clk, f5_11_reg);
        /////////////
        
        assign f6_00 = e_0 ^ eg_0 ^ egh_0 ^ ef_0 ^ d_0 & h_0 ^ d_0 & gh_0 ^ d_0 & fh_0 ^ d_0 & fgh_0 ^ d_0 & eg_0 ^ d_0 & egh_0 ^ d_0 & ef_0 ^ d_0 & efg_0 ^ c_0 ^ c_0 & h_0 ^ c_0 & gh_0 ^ c_0 & fh_0 ^ c_0 & fg_0 ^ c_0 & fgh_0 ^ c_0 & e_0 ^ c_0 & eh_0 ^ c_0 & efh_0 ^ c_0 & efg_0 ^ c_0 & efgh_0 ^ cd_0 & h_0 ^ cd_0 & fh_0 ^ cd_0 & fg_0 ^ cd_0 & egh_0 ^ cd_0 & ef_0 ^ cd_0 & efh_0 ^ cd_0 & efg_0 ^ b_0 ^ b_0 & fh_0 ^ b_0 & fg_0 ^ b_0 & eh_0 ^ b_0 & eg_0 ^ b_0 & egh_0 ^ b_0 & efh_0 ^ b_0 & efg_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & h_0 ^ bd_0 & g_0 ^ bd_0 & f_0 ^ bd_0 & fh_0 ^ bd_0 & e_0 ^ bd_0 & eh_0 ^ bd_0 & eg_0 ^ bd_0 & ef_0 ^ bc_0 & h_0 ^ bc_0 & g_0 ^ bc_0 & ef_0 ^ bc_0 & efh_0 ^ bc_0 & efgh_0 ^ bcd_0 ^ bcd_0 & fg_0 ^ bcd_0 & fgh_0 ^ bcd_0 & eg_0 ^ bcd_0 & egh_0 ^ a_0 & h_0 ^ a_0 & g_0 ^ a_0 & fg_0 ^ a_0 & e_0 ^ a_0 & egh_0 ^ a_0 & ef_0 ^ a_0 & efh_0 ^ a_0 & efgh_0 ^ ad_0 & h_0 ^ ad_0 & g_0 ^ ad_0 & f_0 ^ ad_0 & fg_0 ^ ad_0 & eh_0 ^ ad_0 & eg_0 ^ ad_0 & efg_0 ^ ad_0 & efgh_0 ^ ac_0 ^ ac_0 & h_0 ^ ac_0 & fh_0 ^ ac_0 & e_0 ^ ac_0 & eg_0 ^ ac_0 & ef_0 ^ ac_0 & efg_0 ^ acd_0 & g_0 ^ acd_0 & gh_0 ^ acd_0 & fh_0 ^ acd_0 & fgh_0 ^ acd_0 & eg_0 ^ acd_0 & egh_0 ^ ab_0 & g_0 ^ ab_0 & gh_0 ^ ab_0 & e_0 ^ ab_0 & egh_0 ^ abd_0 & h_0 ^ abd_0 & g_0 ^ abd_0 & fh_0 ^ abd_0 & fgh_0 ^ abd_0 & eh_0 ^ abd_0 & egh_0 ^ abd_0 & ef_0 ^ abc_0 ^ abc_0 & fh_0 ^ abc_0 & fg_0 ^ abc_0 & fgh_0 ^ abc_0 & egh_0 ^ abc_0 & ef_0 ^ abcd_0 ^ abcd_0 & h_0 ^ abcd_0 & g_0 ^ abcd_0 & fgh_0 ^ abcd_0 & e_0 ^ abcd_0 & eg_0 ^ abcd_0 & egh_0 ;
        assign f6_01 = d_0 & h_1 ^ d_0 & gh_1 ^ d_0 & fh_1 ^ d_0 & fgh_1 ^ d_0 & eg_1 ^ d_0 & egh_1 ^ d_0 & ef_1 ^ d_0 & efg_1 ^ c_0 & h_1 ^ c_0 & gh_1 ^ c_0 & fh_1 ^ c_0 & fg_1 ^ c_0 & fgh_1 ^ c_0 & e_1 ^ c_0 & eh_1 ^ c_0 & efh_1 ^ c_0 & efg_1 ^ c_0 & efgh_1 ^ cd_0 & h_1 ^ cd_0 & fh_1 ^ cd_0 & fg_1 ^ cd_0 & egh_1 ^ cd_0 & ef_1 ^ cd_0 & efh_1 ^ cd_0 & efg_1 ^ b_0 & fh_1 ^ b_0 & fg_1 ^ b_0 & eh_1 ^ b_0 & eg_1 ^ b_0 & egh_1 ^ b_0 & efh_1 ^ b_0 & efg_1 ^ b_0 & efgh_1 ^ bd_0 & h_1 ^ bd_0 & g_1 ^ bd_0 & f_1 ^ bd_0 & fh_1 ^ bd_0 & e_1 ^ bd_0 & eh_1 ^ bd_0 & eg_1 ^ bd_0 & ef_1 ^ bc_0 & h_1 ^ bc_0 & g_1 ^ bc_0 & ef_1 ^ bc_0 & efh_1 ^ bc_0 & efgh_1 ^ bcd_0 & fg_1 ^ bcd_0 & fgh_1 ^ bcd_0 & eg_1 ^ bcd_0 & egh_1 ^ a_0 & h_1 ^ a_0 & g_1 ^ a_0 & fg_1 ^ a_0 & e_1 ^ a_0 & egh_1 ^ a_0 & ef_1 ^ a_0 & efh_1 ^ a_0 & efgh_1 ^ ad_0 & h_1 ^ ad_0 & g_1 ^ ad_0 & f_1 ^ ad_0 & fg_1 ^ ad_0 & eh_1 ^ ad_0 & eg_1 ^ ad_0 & efg_1 ^ ad_0 & efgh_1 ^ ac_0 & h_1 ^ ac_0 & fh_1 ^ ac_0 & e_1 ^ ac_0 & eg_1 ^ ac_0 & ef_1 ^ ac_0 & efg_1 ^ acd_0 & g_1 ^ acd_0 & gh_1 ^ acd_0 & fh_1 ^ acd_0 & fgh_1 ^ acd_0 & eg_1 ^ acd_0 & egh_1 ^ ab_0 & g_1 ^ ab_0 & gh_1 ^ ab_0 & e_1 ^ ab_0 & egh_1 ^ abd_0 & h_1 ^ abd_0 & g_1 ^ abd_0 & fh_1 ^ abd_0 & fgh_1 ^ abd_0 & eh_1 ^ abd_0 & egh_1 ^ abd_0 & ef_1 ^ abc_0 & fh_1 ^ abc_0 & fg_1 ^ abc_0 & fgh_1 ^ abc_0 & egh_1 ^ abc_0 & ef_1 ^ abcd_0 & h_1 ^ abcd_0 & g_1 ^ abcd_0 & fgh_1 ^ abcd_0 & e_1 ^ abcd_0 & eg_1 ^ abcd_0 & egh_1 ;
        assign f6_10 = d_1 & h_0 ^ d_1 & gh_0 ^ d_1 & fh_0 ^ d_1 & fgh_0 ^ d_1 & eg_0 ^ d_1 & egh_0 ^ d_1 & ef_0 ^ d_1 & efg_0 ^ c_1 & h_0 ^ c_1 & gh_0 ^ c_1 & fh_0 ^ c_1 & fg_0 ^ c_1 & fgh_0 ^ c_1 & e_0 ^ c_1 & eh_0 ^ c_1 & efh_0 ^ c_1 & efg_0 ^ c_1 & efgh_0 ^ cd_1 & h_0 ^ cd_1 & fh_0 ^ cd_1 & fg_0 ^ cd_1 & egh_0 ^ cd_1 & ef_0 ^ cd_1 & efh_0 ^ cd_1 & efg_0 ^ b_1 & fh_0 ^ b_1 & fg_0 ^ b_1 & eh_0 ^ b_1 & eg_0 ^ b_1 & egh_0 ^ b_1 & efh_0 ^ b_1 & efg_0 ^ b_1 & efgh_0 ^ bd_1 & h_0 ^ bd_1 & g_0 ^ bd_1 & f_0 ^ bd_1 & fh_0 ^ bd_1 & e_0 ^ bd_1 & eh_0 ^ bd_1 & eg_0 ^ bd_1 & ef_0 ^ bc_1 & h_0 ^ bc_1 & g_0 ^ bc_1 & ef_0 ^ bc_1 & efh_0 ^ bc_1 & efgh_0 ^ bcd_1 & fg_0 ^ bcd_1 & fgh_0 ^ bcd_1 & eg_0 ^ bcd_1 & egh_0 ^ a_1 & h_0 ^ a_1 & g_0 ^ a_1 & fg_0 ^ a_1 & e_0 ^ a_1 & egh_0 ^ a_1 & ef_0 ^ a_1 & efh_0 ^ a_1 & efgh_0 ^ ad_1 & h_0 ^ ad_1 & g_0 ^ ad_1 & f_0 ^ ad_1 & fg_0 ^ ad_1 & eh_0 ^ ad_1 & eg_0 ^ ad_1 & efg_0 ^ ad_1 & efgh_0 ^ ac_1 & h_0 ^ ac_1 & fh_0 ^ ac_1 & e_0 ^ ac_1 & eg_0 ^ ac_1 & ef_0 ^ ac_1 & efg_0 ^ acd_1 & g_0 ^ acd_1 & gh_0 ^ acd_1 & fh_0 ^ acd_1 & fgh_0 ^ acd_1 & eg_0 ^ acd_1 & egh_0 ^ ab_1 & g_0 ^ ab_1 & gh_0 ^ ab_1 & e_0 ^ ab_1 & egh_0 ^ abd_1 & h_0 ^ abd_1 & g_0 ^ abd_1 & fh_0 ^ abd_1 & fgh_0 ^ abd_1 & eh_0 ^ abd_1 & egh_0 ^ abd_1 & ef_0 ^ abc_1 & fh_0 ^ abc_1 & fg_0 ^ abc_1 & fgh_0 ^ abc_1 & egh_0 ^ abc_1 & ef_0 ^ abcd_1 & h_0 ^ abcd_1 & g_0 ^ abcd_1 & fgh_0 ^ abcd_1 & e_0 ^ abcd_1 & eg_0 ^ abcd_1 & egh_0 ;
        assign f6_11 = e_1 ^ eg_1 ^ egh_1 ^ ef_1 ^ d_1 & h_1 ^ d_1 & gh_1 ^ d_1 & fh_1 ^ d_1 & fgh_1 ^ d_1 & eg_1 ^ d_1 & egh_1 ^ d_1 & ef_1 ^ d_1 & efg_1 ^ c_1 ^ c_1 & h_1 ^ c_1 & gh_1 ^ c_1 & fh_1 ^ c_1 & fg_1 ^ c_1 & fgh_1 ^ c_1 & e_1 ^ c_1 & eh_1 ^ c_1 & efh_1 ^ c_1 & efg_1 ^ c_1 & efgh_1 ^ cd_1 & h_1 ^ cd_1 & fh_1 ^ cd_1 & fg_1 ^ cd_1 & egh_1 ^ cd_1 & ef_1 ^ cd_1 & efh_1 ^ cd_1 & efg_1 ^ b_1 ^ b_1 & fh_1 ^ b_1 & fg_1 ^ b_1 & eh_1 ^ b_1 & eg_1 ^ b_1 & egh_1 ^ b_1 & efh_1 ^ b_1 & efg_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & h_1 ^ bd_1 & g_1 ^ bd_1 & f_1 ^ bd_1 & fh_1 ^ bd_1 & e_1 ^ bd_1 & eh_1 ^ bd_1 & eg_1 ^ bd_1 & ef_1 ^ bc_1 & h_1 ^ bc_1 & g_1 ^ bc_1 & ef_1 ^ bc_1 & efh_1 ^ bc_1 & efgh_1 ^ bcd_1 ^ bcd_1 & fg_1 ^ bcd_1 & fgh_1 ^ bcd_1 & eg_1 ^ bcd_1 & egh_1 ^ a_1 & h_1 ^ a_1 & g_1 ^ a_1 & fg_1 ^ a_1 & e_1 ^ a_1 & egh_1 ^ a_1 & ef_1 ^ a_1 & efh_1 ^ a_1 & efgh_1 ^ ad_1 & h_1 ^ ad_1 & g_1 ^ ad_1 & f_1 ^ ad_1 & fg_1 ^ ad_1 & eh_1 ^ ad_1 & eg_1 ^ ad_1 & efg_1 ^ ad_1 & efgh_1 ^ ac_1 ^ ac_1 & h_1 ^ ac_1 & fh_1 ^ ac_1 & e_1 ^ ac_1 & eg_1 ^ ac_1 & ef_1 ^ ac_1 & efg_1 ^ acd_1 & g_1 ^ acd_1 & gh_1 ^ acd_1 & fh_1 ^ acd_1 & fgh_1 ^ acd_1 & eg_1 ^ acd_1 & egh_1 ^ ab_1 & g_1 ^ ab_1 & gh_1 ^ ab_1 & e_1 ^ ab_1 & egh_1 ^ abd_1 & h_1 ^ abd_1 & g_1 ^ abd_1 & fh_1 ^ abd_1 & fgh_1 ^ abd_1 & eh_1 ^ abd_1 & egh_1 ^ abd_1 & ef_1 ^ abc_1 ^ abc_1 & fh_1 ^ abc_1 & fg_1 ^ abc_1 & fgh_1 ^ abc_1 & egh_1 ^ abc_1 & ef_1 ^ abcd_1 ^ abcd_1 & h_1 ^ abcd_1 & g_1 ^ abcd_1 & fgh_1 ^ abcd_1 & e_1 ^ abcd_1 & eg_1 ^ abcd_1 & egh_1 ;
        wire f6_00_reg;
        Register # (1) inst_inner_f6_00 (f6_00, clk, f6_00_reg);
        wire f6_01_reg;
        Register # (1) inst_cross_f6_01 (f6_01 ^ r_cross[6], clk, f6_01_reg);
        wire f6_10_reg;
        Register # (1) inst_cross_f6_10 (f6_10 ^ r_cross[6], clk, f6_10_reg);
        wire f6_11_reg;
        Register # (1) inst_inner_f6_11 (f6_11, clk, f6_11_reg);
        //////////////
        
        assign f7_00 = f_0 ^ fh_0 ^ fg_0 ^ efh_0 ^ efg_0 ^ efgh_0 ^ d_0 ^ d_0 & gh_0 ^ d_0 & f_0 ^ d_0 & fgh_0 ^ d_0 & egh_0 ^ d_0 & efg_0 ^ d_0 & efgh_0 ^ c_0 ^ c_0 & gh_0 ^ c_0 & fh_0 ^ c_0 & fgh_0 ^ c_0 & e_0 ^ c_0 & eh_0 ^ c_0 & eg_0 ^ c_0 & ef_0 ^ c_0 & efh_0 ^ c_0 & efg_0 ^ cd_0 & h_0 ^ cd_0 & fg_0 ^ cd_0 & e_0 ^ cd_0 & egh_0 ^ cd_0 & efh_0 ^ b_0 & h_0 ^ b_0 & gh_0 ^ b_0 & f_0 ^ b_0 & fg_0 ^ b_0 & eh_0 ^ b_0 & eg_0 ^ b_0 & egh_0 ^ b_0 & efh_0 ^ b_0 & efgh_0 ^ bd_0 ^ bd_0 & f_0 ^ bd_0 & fh_0 ^ bd_0 & fg_0 ^ bd_0 & fgh_0 ^ bd_0 & eh_0 ^ bd_0 & efh_0 ^ bc_0 & h_0 ^ bc_0 & f_0 ^ bc_0 & eh_0 ^ bc_0 & efg_0 ^ bcd_0 ^ bcd_0 & gh_0 ^ bcd_0 & fg_0 ^ bcd_0 & e_0 ^ bcd_0 & eh_0 ^ bcd_0 & ef_0 ^ bcd_0 & efh_0 ^ a_0 ^ a_0 & h_0 ^ a_0 & g_0 ^ a_0 & fh_0 ^ a_0 & fgh_0 ^ a_0 & eh_0 ^ a_0 & efh_0 ^ a_0 & efg_0 ^ ad_0 & g_0 ^ ad_0 & gh_0 ^ ad_0 & fh_0 ^ ad_0 & eh_0 ^ ad_0 & eg_0 ^ ad_0 & egh_0 ^ ad_0 & ef_0 ^ ad_0 & efh_0 ^ ac_0 ^ ac_0 & fgh_0 ^ ac_0 & e_0 ^ ac_0 & eh_0 ^ acd_0 ^ acd_0 & g_0 ^ acd_0 & gh_0 ^ acd_0 & fgh_0 ^ acd_0 & egh_0 ^ acd_0 & efh_0 ^ ab_0 & h_0 ^ ab_0 & f_0 ^ ab_0 & fgh_0 ^ ab_0 & eh_0 ^ ab_0 & eg_0 ^ ab_0 & efgh_0 ^ abd_0 ^ abd_0 & h_0 ^ abd_0 & g_0 ^ abd_0 & f_0 ^ abd_0 & fg_0 ^ abd_0 & eh_0 ^ abd_0 & egh_0 ^ abd_0 & efh_0 ^ abc_0 & g_0 ^ abc_0 & gh_0 ^ abc_0 & f_0 ^ abc_0 & fg_0 ^ abc_0 & eh_0 ^ abc_0 & eg_0 ^ abc_0 & egh_0 ^ abc_0 & efh_0 ^ abcd_0 ^ abcd_0 & g_0 ^ abcd_0 & fh_0 ^ abcd_0 & e_0 ^ abcd_0 & eg_0 ^ abcd_0 & egh_0 ^ abcd_0 & efh_0 ;
        assign f7_01 = d_0 & gh_1 ^ d_0 & f_1 ^ d_0 & fgh_1 ^ d_0 & egh_1 ^ d_0 & efg_1 ^ d_0 & efgh_1 ^ c_0 & gh_1 ^ c_0 & fh_1 ^ c_0 & fgh_1 ^ c_0 & e_1 ^ c_0 & eh_1 ^ c_0 & eg_1 ^ c_0 & ef_1 ^ c_0 & efh_1 ^ c_0 & efg_1 ^ cd_0 & h_1 ^ cd_0 & fg_1 ^ cd_0 & e_1 ^ cd_0 & egh_1 ^ cd_0 & efh_1 ^ b_0 & h_1 ^ b_0 & gh_1 ^ b_0 & f_1 ^ b_0 & fg_1 ^ b_0 & eh_1 ^ b_0 & eg_1 ^ b_0 & egh_1 ^ b_0 & efh_1 ^ b_0 & efgh_1 ^ bd_0 & f_1 ^ bd_0 & fh_1 ^ bd_0 & fg_1 ^ bd_0 & fgh_1 ^ bd_0 & eh_1 ^ bd_0 & efh_1 ^ bc_0 & h_1 ^ bc_0 & f_1 ^ bc_0 & eh_1 ^ bc_0 & efg_1 ^ bcd_0 & gh_1 ^ bcd_0 & fg_1 ^ bcd_0 & e_1 ^ bcd_0 & eh_1 ^ bcd_0 & ef_1 ^ bcd_0 & efh_1 ^ a_0 & h_1 ^ a_0 & g_1 ^ a_0 & fh_1 ^ a_0 & fgh_1 ^ a_0 & eh_1 ^ a_0 & efh_1 ^ a_0 & efg_1 ^ ad_0 & g_1 ^ ad_0 & gh_1 ^ ad_0 & fh_1 ^ ad_0 & eh_1 ^ ad_0 & eg_1 ^ ad_0 & egh_1 ^ ad_0 & ef_1 ^ ad_0 & efh_1 ^ ac_0 & fgh_1 ^ ac_0 & e_1 ^ ac_0 & eh_1 ^ acd_0 & g_1 ^ acd_0 & gh_1 ^ acd_0 & fgh_1 ^ acd_0 & egh_1 ^ acd_0 & efh_1 ^ ab_0 & h_1 ^ ab_0 & f_1 ^ ab_0 & fgh_1 ^ ab_0 & eh_1 ^ ab_0 & eg_1 ^ ab_0 & efgh_1 ^ abd_0 & h_1 ^ abd_0 & g_1 ^ abd_0 & f_1 ^ abd_0 & fg_1 ^ abd_0 & eh_1 ^ abd_0 & egh_1 ^ abd_0 & efh_1 ^ abc_0 & g_1 ^ abc_0 & gh_1 ^ abc_0 & f_1 ^ abc_0 & fg_1 ^ abc_0 & eh_1 ^ abc_0 & eg_1 ^ abc_0 & egh_1 ^ abc_0 & efh_1 ^ abcd_0 & g_1 ^ abcd_0 & fh_1 ^ abcd_0 & e_1 ^ abcd_0 & eg_1 ^ abcd_0 & egh_1 ^ abcd_0 & efh_1 ;
        assign f7_10 = d_1 & gh_0 ^ d_1 & f_0 ^ d_1 & fgh_0 ^ d_1 & egh_0 ^ d_1 & efg_0 ^ d_1 & efgh_0 ^ c_1 & gh_0 ^ c_1 & fh_0 ^ c_1 & fgh_0 ^ c_1 & e_0 ^ c_1 & eh_0 ^ c_1 & eg_0 ^ c_1 & ef_0 ^ c_1 & efh_0 ^ c_1 & efg_0 ^ cd_1 & h_0 ^ cd_1 & fg_0 ^ cd_1 & e_0 ^ cd_1 & egh_0 ^ cd_1 & efh_0 ^ b_1 & h_0 ^ b_1 & gh_0 ^ b_1 & f_0 ^ b_1 & fg_0 ^ b_1 & eh_0 ^ b_1 & eg_0 ^ b_1 & egh_0 ^ b_1 & efh_0 ^ b_1 & efgh_0 ^ bd_1 & f_0 ^ bd_1 & fh_0 ^ bd_1 & fg_0 ^ bd_1 & fgh_0 ^ bd_1 & eh_0 ^ bd_1 & efh_0 ^ bc_1 & h_0 ^ bc_1 & f_0 ^ bc_1 & eh_0 ^ bc_1 & efg_0 ^ bcd_1 & gh_0 ^ bcd_1 & fg_0 ^ bcd_1 & e_0 ^ bcd_1 & eh_0 ^ bcd_1 & ef_0 ^ bcd_1 & efh_0 ^ a_1 & h_0 ^ a_1 & g_0 ^ a_1 & fh_0 ^ a_1 & fgh_0 ^ a_1 & eh_0 ^ a_1 & efh_0 ^ a_1 & efg_0 ^ ad_1 & g_0 ^ ad_1 & gh_0 ^ ad_1 & fh_0 ^ ad_1 & eh_0 ^ ad_1 & eg_0 ^ ad_1 & egh_0 ^ ad_1 & ef_0 ^ ad_1 & efh_0 ^ ac_1 & fgh_0 ^ ac_1 & e_0 ^ ac_1 & eh_0 ^ acd_1 & g_0 ^ acd_1 & gh_0 ^ acd_1 & fgh_0 ^ acd_1 & egh_0 ^ acd_1 & efh_0 ^ ab_1 & h_0 ^ ab_1 & f_0 ^ ab_1 & fgh_0 ^ ab_1 & eh_0 ^ ab_1 & eg_0 ^ ab_1 & efgh_0 ^ abd_1 & h_0 ^ abd_1 & g_0 ^ abd_1 & f_0 ^ abd_1 & fg_0 ^ abd_1 & eh_0 ^ abd_1 & egh_0 ^ abd_1 & efh_0 ^ abc_1 & g_0 ^ abc_1 & gh_0 ^ abc_1 & f_0 ^ abc_1 & fg_0 ^ abc_1 & eh_0 ^ abc_1 & eg_0 ^ abc_1 & egh_0 ^ abc_1 & efh_0 ^ abcd_1 & g_0 ^ abcd_1 & fh_0 ^ abcd_1 & e_0 ^ abcd_1 & eg_0 ^ abcd_1 & egh_0 ^ abcd_1 & efh_0 ;
        assign f7_11 = f_1 ^ fh_1 ^ fg_1 ^ efh_1 ^ efg_1 ^ efgh_1 ^ d_1 ^ d_1 & gh_1 ^ d_1 & f_1 ^ d_1 & fgh_1 ^ d_1 & egh_1 ^ d_1 & efg_1 ^ d_1 & efgh_1 ^ c_1 ^ c_1 & gh_1 ^ c_1 & fh_1 ^ c_1 & fgh_1 ^ c_1 & e_1 ^ c_1 & eh_1 ^ c_1 & eg_1 ^ c_1 & ef_1 ^ c_1 & efh_1 ^ c_1 & efg_1 ^ cd_1 & h_1 ^ cd_1 & fg_1 ^ cd_1 & e_1 ^ cd_1 & egh_1 ^ cd_1 & efh_1 ^ b_1 & h_1 ^ b_1 & gh_1 ^ b_1 & f_1 ^ b_1 & fg_1 ^ b_1 & eh_1 ^ b_1 & eg_1 ^ b_1 & egh_1 ^ b_1 & efh_1 ^ b_1 & efgh_1 ^ bd_1 ^ bd_1 & f_1 ^ bd_1 & fh_1 ^ bd_1 & fg_1 ^ bd_1 & fgh_1 ^ bd_1 & eh_1 ^ bd_1 & efh_1 ^ bc_1 & h_1 ^ bc_1 & f_1 ^ bc_1 & eh_1 ^ bc_1 & efg_1 ^ bcd_1 ^ bcd_1 & gh_1 ^ bcd_1 & fg_1 ^ bcd_1 & e_1 ^ bcd_1 & eh_1 ^ bcd_1 & ef_1 ^ bcd_1 & efh_1 ^ a_1 ^ a_1 & h_1 ^ a_1 & g_1 ^ a_1 & fh_1 ^ a_1 & fgh_1 ^ a_1 & eh_1 ^ a_1 & efh_1 ^ a_1 & efg_1 ^ ad_1 & g_1 ^ ad_1 & gh_1 ^ ad_1 & fh_1 ^ ad_1 & eh_1 ^ ad_1 & eg_1 ^ ad_1 & egh_1 ^ ad_1 & ef_1 ^ ad_1 & efh_1 ^ ac_1 ^ ac_1 & fgh_1 ^ ac_1 & e_1 ^ ac_1 & eh_1 ^ acd_1 ^ acd_1 & g_1 ^ acd_1 & gh_1 ^ acd_1 & fgh_1 ^ acd_1 & egh_1 ^ acd_1 & efh_1 ^ ab_1 & h_1 ^ ab_1 & f_1 ^ ab_1 & fgh_1 ^ ab_1 & eh_1 ^ ab_1 & eg_1 ^ ab_1 & efgh_1 ^ abd_1 ^ abd_1 & h_1 ^ abd_1 & g_1 ^ abd_1 & f_1 ^ abd_1 & fg_1 ^ abd_1 & eh_1 ^ abd_1 & egh_1 ^ abd_1 & efh_1 ^ abc_1 & g_1 ^ abc_1 & gh_1 ^ abc_1 & f_1 ^ abc_1 & fg_1 ^ abc_1 & eh_1 ^ abc_1 & eg_1 ^ abc_1 & egh_1 ^ abc_1 & efh_1 ^ abcd_1 ^ abcd_1 & g_1 ^ abcd_1 & fh_1 ^ abcd_1 & e_1 ^ abcd_1 & eg_1 ^ abcd_1 & egh_1 ^ abcd_1 & efh_1 ;
        wire f7_00_reg;
        Register # (1) inst_inner_f7_00 (f7_00, clk, f7_00_reg);
        wire f7_01_reg;
        Register # (1) inst_cross_f7_01 (f7_01 ^ r_cross[7], clk, f7_01_reg);
        wire f7_10_reg;
        Register # (1) inst_cross_f7_10 (f7_10 ^ r_cross[7], clk, f7_10_reg);
        wire f7_11_reg;
        Register # (1) inst_inner_f7_11 (f7_11, clk, f7_11_reg);
        //////////////
        
        
        assign F0[0] = f0_00_reg ^ f0_01_reg;
        assign F1[0] = f0_10_reg ^ f0_11_reg ^ 1'b1;
        
        assign F0[1] = f1_00_reg ^ f1_01_reg;
        assign F1[1] = f1_10_reg ^ f1_11_reg ^ 1'b1;
        
        assign F0[2] = f2_00_reg ^ f2_01_reg;
        assign F1[2] = f2_10_reg ^ f2_11_reg;
        
        assign F0[3] = f3_00_reg ^ f3_01_reg;
        assign F1[3] = f3_10_reg ^ f3_11_reg;
        
        assign F0[4] = f4_00_reg ^ f4_01_reg;
        assign F1[4] = f4_10_reg ^ f4_11_reg;
        
        assign F0[5] = f5_00_reg ^ f5_01_reg;
        assign F1[5] = f5_10_reg ^ f5_11_reg ^ 1'b1;
        
        assign F0[6] = f6_00_reg ^ f6_01_reg;
        assign F1[6] = f6_10_reg ^ f6_11_reg ^ 1'b1;
        
        assign F0[7] = f7_00_reg ^ f7_01_reg;
        assign F1[7] = f7_10_reg ^ f7_11_reg;
        
endmodule
